module assertion_gen();

`define ADC0EXTMUXSEL0_IN 0
`define ADC0EXTMUXSEL0_OE 0
`define ADC0EXTMUXSEL0_OUT 0
`define ADC0EXTMUXSEL1_IN 0
`define ADC0EXTMUXSEL1_OE 0
`define ADC0EXTMUXSEL1_OUT 0
`define ADC0EXTMUXSEL2_IN 0
`define ADC0EXTMUXSEL2_OE 0
`define ADC0EXTMUXSEL2_OUT 0
`define ADC0EXTMUXSEL3_IN 0
`define ADC0EXTMUXSEL3_OE 0
`define ADC0EXTMUXSEL3_OUT 0
`define ADC1EXTMUXSEL0_IN 0
`define ADC1EXTMUXSEL0_OE 0
`define ADC1EXTMUXSEL0_OUT 0
`define ADC1EXTMUXSEL1_IN 0
`define ADC1EXTMUXSEL1_OE 0
`define ADC1EXTMUXSEL1_OUT 0
`define ADC1EXTMUXSEL2_IN 0
`define ADC1EXTMUXSEL2_OE 0
`define ADC1EXTMUXSEL2_OUT 0
`define ADC1EXTMUXSEL3_IN 0
`define ADC1EXTMUXSEL3_OE 0
`define ADC1EXTMUXSEL3_OUT 0
`define ADC2EXTMUXSEL0_IN 0
`define ADC2EXTMUXSEL0_OE 0
`define ADC2EXTMUXSEL0_OUT 0
`define ADC2EXTMUXSEL1_IN 0
`define ADC2EXTMUXSEL1_OE 0
`define ADC2EXTMUXSEL1_OUT 0
`define ADC2EXTMUXSEL2_IN 0
`define ADC2EXTMUXSEL2_OE 0
`define ADC2EXTMUXSEL2_OUT 0
`define ADC2EXTMUXSEL3_IN 0
`define ADC2EXTMUXSEL3_OE 0
`define ADC2EXTMUXSEL3_OUT 0
`define ADC3EXTMUXSEL0_IN 0
`define ADC3EXTMUXSEL0_OE 0
`define ADC3EXTMUXSEL0_OUT 0
`define ADC3EXTMUXSEL1_IN 0
`define ADC3EXTMUXSEL1_OE 0
`define ADC3EXTMUXSEL1_OUT 0
`define ADC3EXTMUXSEL2_IN 0
`define ADC3EXTMUXSEL2_OE 0
`define ADC3EXTMUXSEL2_OUT 0
`define ADC3EXTMUXSEL3_IN 0
`define ADC3EXTMUXSEL3_OE 0
`define ADC3EXTMUXSEL3_OUT 0
`define ADC4EXTMUXSEL0_IN 0
`define ADC4EXTMUXSEL0_OE 0
`define ADC4EXTMUXSEL0_OUT 0
`define ADC4EXTMUXSEL1_IN 0
`define ADC4EXTMUXSEL1_OE 0
`define ADC4EXTMUXSEL1_OUT 0
`define ADC4EXTMUXSEL2_IN 0
`define ADC4EXTMUXSEL2_OE 0
`define ADC4EXTMUXSEL2_OUT 0
`define ADC4EXTMUXSEL3_IN 0
`define ADC4EXTMUXSEL3_OE 0
`define ADC4EXTMUXSEL3_OUT 0
`define ADC5EXTMUXSEL0_IN 0
`define ADC5EXTMUXSEL0_OE 0
`define ADC5EXTMUXSEL0_OUT 0
`define ADC5EXTMUXSEL1_IN 0
`define ADC5EXTMUXSEL1_OE 0
`define ADC5EXTMUXSEL1_OUT 0
`define ADC5EXTMUXSEL2_IN 0
`define ADC5EXTMUXSEL2_OE 0
`define ADC5EXTMUXSEL2_OUT 0
`define ADC5EXTMUXSEL3_IN 0
`define ADC5EXTMUXSEL3_OE 0
`define ADC5EXTMUXSEL3_OUT 0
`define ADC6EXTMUXSEL0_IN 0
`define ADC6EXTMUXSEL0_OE 0
`define ADC6EXTMUXSEL0_OUT 0
`define ADC6EXTMUXSEL1_IN 0
`define ADC6EXTMUXSEL1_OE 0
`define ADC6EXTMUXSEL1_OUT 0
`define ADC6EXTMUXSEL2_IN 0
`define ADC6EXTMUXSEL2_OE 0
`define ADC6EXTMUXSEL2_OUT 0
`define ADC6EXTMUXSEL3_IN 0
`define ADC6EXTMUXSEL3_OE 0
`define ADC6EXTMUXSEL3_OUT 0
`define ADC7EXTMUXSEL0_IN 0
`define ADC7EXTMUXSEL0_OE 0
`define ADC7EXTMUXSEL0_OUT 0
`define ADC7EXTMUXSEL1_IN 0
`define ADC7EXTMUXSEL1_OE 0
`define ADC7EXTMUXSEL1_OUT 0
`define ADC7EXTMUXSEL2_IN 0
`define ADC7EXTMUXSEL2_OE 0
`define ADC7EXTMUXSEL2_OUT 0
`define ADC7EXTMUXSEL3_IN 0
`define ADC7EXTMUXSEL3_OE 0
`define ADC7EXTMUXSEL3_OUT 0
`define ADCSOC0_IN 0
`define ADCSOC0_OE 0
`define ADCSOC0_OUT 0
`define ADCSOC1_IN 0
`define ADCSOC1_OE 0
`define ADCSOC1_OUT 0
`define CAN0RX_IN 0
`define CAN0RX_OE 0
`define CAN0RX_OUT 0
`define CAN0TX_IN 0
`define CAN0TX_OE 0
`define CAN0TX_OUT 0
`define CAN10RX_IN 0
`define CAN10RX_OE 0
`define CAN10RX_OUT 0
`define CAN10TX_IN 0
`define CAN10TX_OE 0
`define CAN10TX_OUT 0
`define CAN11RX_IN 0
`define CAN11RX_OE 0
`define CAN11RX_OUT 0
`define CAN11TX_IN 0
`define CAN11TX_OE 0
`define CAN11TX_OUT 0
`define CAN1RX_IN 0
`define CAN1RX_OE 0
`define CAN1RX_OUT 0
`define CAN1TX_IN 0
`define CAN1TX_OE 0
`define CAN1TX_OUT 0
`define CAN2RX_IN 0
`define CAN2RX_OE 0
`define CAN2RX_OUT 0
`define CAN2TX_IN 0
`define CAN2TX_OE 0
`define CAN2TX_OUT 0
`define CAN3RX_IN 0
`define CAN3RX_OE 0
`define CAN3RX_OUT 0
`define CAN3TX_IN 0
`define CAN3TX_OE 0
`define CAN3TX_OUT 0
`define CAN4RX_IN 0
`define CAN4RX_OE 0
`define CAN4RX_OUT 0
`define CAN4TX_IN 0
`define CAN4TX_OE 0
`define CAN4TX_OUT 0
`define CAN5RX_IN 0
`define CAN5RX_OE 0
`define CAN5RX_OUT 0
`define CAN5TX_IN 0
`define CAN5TX_OE 0
`define CAN5TX_OUT 0
`define CAN6RX_IN 0
`define CAN6RX_OE 0
`define CAN6RX_OUT 0
`define CAN6TX_IN 0
`define CAN6TX_OE 0
`define CAN6TX_OUT 0
`define CAN7RX_IN 0
`define CAN7RX_OE 0
`define CAN7RX_OUT 0
`define CAN7TX_IN 0
`define CAN7TX_OE 0
`define CAN7TX_OUT 0
`define CAN8RX_IN 0
`define CAN8RX_OE 0
`define CAN8RX_OUT 0
`define CAN8TX_IN 0
`define CAN8TX_OE 0
`define CAN8TX_OUT 0
`define CAN9RX_IN 0
`define CAN9RX_OE 0
`define CAN9RX_OUT 0
`define CAN9TX_IN 0
`define CAN9TX_OE 0
`define CAN9TX_OUT 0
`define CLKOUT1_IN 0
`define CLKOUT1_OE 0
`define CLKOUT1_OUT 0
`define CLKOUT2_IN 0
`define CLKOUT2_OE 0
`define CLKOUT2_OUT 0
`define DP0_0 0
`define DP0_0_GPIO_OUTPUT_ENABLE 0
`define DP0_0_INFUNC_EN 0
`define DP0_0_OUTFUNC_SEL 0
`define DP0_0_PINCTRL_0_IE 0
`define DP0_0_PINCTRL_0_OD 0
`define DP0_0_PULLEN 0
`define DP0_0_PULLSEL 0
`define DP0_0_pad_y 0
`define DP0_1 0
`define DP0_10 0
`define DP0_10_GPIO_OUTPUT_ENABLE 0
`define DP0_10_INFUNC_EN 0
`define DP0_10_OUTFUNC_SEL 0
`define DP0_10_PINCTRL_0_IE 0
`define DP0_10_PINCTRL_0_OD 0
`define DP0_10_PULLEN 0
`define DP0_10_PULLSEL 0
`define DP0_10_pad_y 0
`define DP0_11 0
`define DP0_11_GPIO_OUTPUT_ENABLE 0
`define DP0_11_INFUNC_EN 0
`define DP0_11_OUTFUNC_SEL 0
`define DP0_11_PINCTRL_0_IE 0
`define DP0_11_PINCTRL_0_OD 0
`define DP0_11_PULLEN 0
`define DP0_11_PULLSEL 0
`define DP0_11_pad_y 0
`define DP0_12 0
`define DP0_12_GPIO_OUTPUT_ENABLE 0
`define DP0_12_INFUNC_EN 0
`define DP0_12_OUTFUNC_SEL 0
`define DP0_12_PINCTRL_0_IE 0
`define DP0_12_PINCTRL_0_OD 0
`define DP0_12_PULLEN 0
`define DP0_12_PULLSEL 0
`define DP0_12_pad_y 0
`define DP0_13 0
`define DP0_13_GPIO_OUTPUT_ENABLE 0
`define DP0_13_INFUNC_EN 0
`define DP0_13_OUTFUNC_SEL 0
`define DP0_13_PINCTRL_0_IE 0
`define DP0_13_PINCTRL_0_OD 0
`define DP0_13_PULLEN 0
`define DP0_13_PULLSEL 0
`define DP0_13_pad_y 0
`define DP0_14 0
`define DP0_14_GPIO_OUTPUT_ENABLE 0
`define DP0_14_INFUNC_EN 0
`define DP0_14_OUTFUNC_SEL 0
`define DP0_14_PINCTRL_0_IE 0
`define DP0_14_PINCTRL_0_OD 0
`define DP0_14_PULLEN 0
`define DP0_14_PULLSEL 0
`define DP0_14_pad_y 0
`define DP0_15 0
`define DP0_15_GPIO_OUTPUT_ENABLE 0
`define DP0_15_INFUNC_EN 0
`define DP0_15_OUTFUNC_SEL 0
`define DP0_15_PINCTRL_0_IE 0
`define DP0_15_PINCTRL_0_OD 0
`define DP0_15_PULLEN 0
`define DP0_15_PULLSEL 0
`define DP0_15_pad_y 0
`define DP0_16 0
`define DP0_16_GPIO_OUTPUT_ENABLE 0
`define DP0_16_INFUNC_EN 0
`define DP0_16_OUTFUNC_SEL 0
`define DP0_16_PINCTRL_0_IE 0
`define DP0_16_PINCTRL_0_OD 0
`define DP0_16_PULLEN 0
`define DP0_16_PULLSEL 0
`define DP0_16_pad_y 0
`define DP0_17 0
`define DP0_17_GPIO_OUTPUT_ENABLE 0
`define DP0_17_INFUNC_EN 0
`define DP0_17_OUTFUNC_SEL 0
`define DP0_17_PINCTRL_0_IE 0
`define DP0_17_PINCTRL_0_OD 0
`define DP0_17_PULLEN 0
`define DP0_17_PULLSEL 0
`define DP0_17_pad_y 0
`define DP0_18 0
`define DP0_18_GPIO_OUTPUT_ENABLE 0
`define DP0_18_INFUNC_EN 0
`define DP0_18_OUTFUNC_SEL 0
`define DP0_18_PINCTRL_0_IE 0
`define DP0_18_PINCTRL_0_OD 0
`define DP0_18_PULLEN 0
`define DP0_18_PULLSEL 0
`define DP0_18_pad_y 0
`define DP0_19 0
`define DP0_19_GPIO_OUTPUT_ENABLE 0
`define DP0_19_INFUNC_EN 0
`define DP0_19_OUTFUNC_SEL 0
`define DP0_19_PINCTRL_0_IE 0
`define DP0_19_PINCTRL_0_OD 0
`define DP0_19_PULLEN 0
`define DP0_19_PULLSEL 0
`define DP0_19_pad_y 0
`define DP0_1_GPIO_OUTPUT_ENABLE 0
`define DP0_1_INFUNC_EN 0
`define DP0_1_OUTFUNC_SEL 0
`define DP0_1_PINCTRL_0_IE 0
`define DP0_1_PINCTRL_0_OD 0
`define DP0_1_PULLEN 0
`define DP0_1_PULLSEL 0
`define DP0_1_pad_y 0
`define DP0_2 0
`define DP0_20 0
`define DP0_20_GPIO_OUTPUT_ENABLE 0
`define DP0_20_INFUNC_EN 0
`define DP0_20_OUTFUNC_SEL 0
`define DP0_20_PINCTRL_0_IE 0
`define DP0_20_PINCTRL_0_OD 0
`define DP0_20_PULLEN 0
`define DP0_20_PULLSEL 0
`define DP0_20_pad_y 0
`define DP0_21 0
`define DP0_21_GPIO_OUTPUT_ENABLE 0
`define DP0_21_INFUNC_EN 0
`define DP0_21_OUTFUNC_SEL 0
`define DP0_21_PINCTRL_0_IE 0
`define DP0_21_PINCTRL_0_OD 0
`define DP0_21_PULLEN 0
`define DP0_21_PULLSEL 0
`define DP0_21_pad_y 0
`define DP0_22 0
`define DP0_22_GPIO_OUTPUT_ENABLE 0
`define DP0_22_INFUNC_EN 0
`define DP0_22_OUTFUNC_SEL 0
`define DP0_22_PINCTRL_0_IE 0
`define DP0_22_PINCTRL_0_OD 0
`define DP0_22_PULLEN 0
`define DP0_22_PULLSEL 0
`define DP0_22_pad_y 0
`define DP0_23 0
`define DP0_23_GPIO_OUTPUT_ENABLE 0
`define DP0_23_INFUNC_EN 0
`define DP0_23_OUTFUNC_SEL 0
`define DP0_23_PINCTRL_0_IE 0
`define DP0_23_PINCTRL_0_OD 0
`define DP0_23_PULLEN 0
`define DP0_23_PULLSEL 0
`define DP0_23_pad_y 0
`define DP0_24 0
`define DP0_24_GPIO_OUTPUT_ENABLE 0
`define DP0_24_INFUNC_EN 0
`define DP0_24_OUTFUNC_SEL 0
`define DP0_24_PINCTRL_0_IE 0
`define DP0_24_PINCTRL_0_OD 0
`define DP0_24_PULLEN 0
`define DP0_24_PULLSEL 0
`define DP0_24_pad_y 0
`define DP0_25 0
`define DP0_25_GPIO_OUTPUT_ENABLE 0
`define DP0_25_INFUNC_EN 0
`define DP0_25_OUTFUNC_SEL 0
`define DP0_25_PINCTRL_0_IE 0
`define DP0_25_PINCTRL_0_OD 0
`define DP0_25_PULLEN 0
`define DP0_25_PULLSEL 0
`define DP0_25_pad_y 0
`define DP0_26 0
`define DP0_26_GPIO_OUTPUT_ENABLE 0
`define DP0_26_INFUNC_EN 0
`define DP0_26_OUTFUNC_SEL 0
`define DP0_26_PINCTRL_0_IE 0
`define DP0_26_PINCTRL_0_OD 0
`define DP0_26_PULLEN 0
`define DP0_26_PULLSEL 0
`define DP0_26_pad_y 0
`define DP0_27 0
`define DP0_27_GPIO_OUTPUT_ENABLE 0
`define DP0_27_INFUNC_EN 0
`define DP0_27_OUTFUNC_SEL 0
`define DP0_27_PINCTRL_0_IE 0
`define DP0_27_PINCTRL_0_OD 0
`define DP0_27_PULLEN 0
`define DP0_27_PULLSEL 0
`define DP0_27_pad_y 0
`define DP0_28 0
`define DP0_28_GPIO_OUTPUT_ENABLE 0
`define DP0_28_INFUNC_EN 0
`define DP0_28_OUTFUNC_SEL 0
`define DP0_28_PINCTRL_0_IE 0
`define DP0_28_PINCTRL_0_OD 0
`define DP0_28_PULLEN 0
`define DP0_28_PULLSEL 0
`define DP0_28_pad_y 0
`define DP0_29 0
`define DP0_29_GPIO_OUTPUT_ENABLE 0
`define DP0_29_INFUNC_EN 0
`define DP0_29_OUTFUNC_SEL 0
`define DP0_29_PINCTRL_0_IE 0
`define DP0_29_PINCTRL_0_OD 0
`define DP0_29_PULLEN 0
`define DP0_29_PULLSEL 0
`define DP0_29_pad_y 0
`define DP0_2_GPIO_OUTPUT_ENABLE 0
`define DP0_2_INFUNC_EN 0
`define DP0_2_OUTFUNC_SEL 0
`define DP0_2_PINCTRL_0_IE 0
`define DP0_2_PINCTRL_0_OD 0
`define DP0_2_PULLEN 0
`define DP0_2_PULLSEL 0
`define DP0_2_pad_y 0
`define DP0_3 0
`define DP0_30 0
`define DP0_30_GPIO_OUTPUT_ENABLE 0
`define DP0_30_INFUNC_EN 0
`define DP0_30_OUTFUNC_SEL 0
`define DP0_30_PINCTRL_0_IE 0
`define DP0_30_PINCTRL_0_OD 0
`define DP0_30_PULLEN 0
`define DP0_30_PULLSEL 0
`define DP0_30_pad_y 0
`define DP0_31 0
`define DP0_31_GPIO_OUTPUT_ENABLE 0
`define DP0_31_INFUNC_EN 0
`define DP0_31_OUTFUNC_SEL 0
`define DP0_31_PINCTRL_0_IE 0
`define DP0_31_PINCTRL_0_OD 0
`define DP0_31_PULLEN 0
`define DP0_31_PULLSEL 0
`define DP0_31_pad_y 0
`define DP0_3_GPIO_OUTPUT_ENABLE 0
`define DP0_3_INFUNC_EN 0
`define DP0_3_OUTFUNC_SEL 0
`define DP0_3_PINCTRL_0_IE 0
`define DP0_3_PINCTRL_0_OD 0
`define DP0_3_PULLEN 0
`define DP0_3_PULLSEL 0
`define DP0_3_pad_y 0
`define DP0_4 0
`define DP0_4_GPIO_OUTPUT_ENABLE 0
`define DP0_4_INFUNC_EN 0
`define DP0_4_OUTFUNC_SEL 0
`define DP0_4_PINCTRL_0_IE 0
`define DP0_4_PINCTRL_0_OD 0
`define DP0_4_PULLEN 0
`define DP0_4_PULLSEL 0
`define DP0_4_pad_y 0
`define DP0_5 0
`define DP0_5_GPIO_OUTPUT_ENABLE 0
`define DP0_5_INFUNC_EN 0
`define DP0_5_OUTFUNC_SEL 0
`define DP0_5_PINCTRL_0_IE 0
`define DP0_5_PINCTRL_0_OD 0
`define DP0_5_PULLEN 0
`define DP0_5_PULLSEL 0
`define DP0_5_pad_y 0
`define DP0_6 0
`define DP0_6_GPIO_OUTPUT_ENABLE 0
`define DP0_6_INFUNC_EN 0
`define DP0_6_OUTFUNC_SEL 0
`define DP0_6_PINCTRL_0_IE 0
`define DP0_6_PINCTRL_0_OD 0
`define DP0_6_PULLEN 0
`define DP0_6_PULLSEL 0
`define DP0_6_pad_y 0
`define DP0_7 0
`define DP0_7_GPIO_OUTPUT_ENABLE 0
`define DP0_7_INFUNC_EN 0
`define DP0_7_OUTFUNC_SEL 0
`define DP0_7_PINCTRL_0_IE 0
`define DP0_7_PINCTRL_0_OD 0
`define DP0_7_PULLEN 0
`define DP0_7_PULLSEL 0
`define DP0_7_pad_y 0
`define DP0_8 0
`define DP0_8_GPIO_OUTPUT_ENABLE 0
`define DP0_8_INFUNC_EN 0
`define DP0_8_OUTFUNC_SEL 0
`define DP0_8_PINCTRL_0_IE 0
`define DP0_8_PINCTRL_0_OD 0
`define DP0_8_PULLEN 0
`define DP0_8_PULLSEL 0
`define DP0_8_pad_y 0
`define DP0_9 0
`define DP0_9_GPIO_OUTPUT_ENABLE 0
`define DP0_9_INFUNC_EN 0
`define DP0_9_OUTFUNC_SEL 0
`define DP0_9_PINCTRL_0_IE 0
`define DP0_9_PINCTRL_0_OD 0
`define DP0_9_PULLEN 0
`define DP0_9_PULLSEL 0
`define DP0_9_pad_y 0
`define DP1_0 0
`define DP1_0_GPIO_OUTPUT_ENABLE 0
`define DP1_0_INFUNC_EN 0
`define DP1_0_OUTFUNC_SEL 0
`define DP1_0_PINCTRL_0_IE 0
`define DP1_0_PINCTRL_0_OD 0
`define DP1_0_PULLEN 0
`define DP1_0_PULLSEL 0
`define DP1_0_pad_y 0
`define DP1_1 0
`define DP1_10 0
`define DP1_10_GPIO_OUTPUT_ENABLE 0
`define DP1_10_INFUNC_EN 0
`define DP1_10_OUTFUNC_SEL 0
`define DP1_10_PINCTRL_0_IE 0
`define DP1_10_PINCTRL_0_OD 0
`define DP1_10_PULLEN 0
`define DP1_10_PULLSEL 0
`define DP1_10_pad_y 0
`define DP1_11 0
`define DP1_11_GPIO_OUTPUT_ENABLE 0
`define DP1_11_INFUNC_EN 0
`define DP1_11_OUTFUNC_SEL 0
`define DP1_11_PINCTRL_0_IE 0
`define DP1_11_PINCTRL_0_OD 0
`define DP1_11_PULLEN 0
`define DP1_11_PULLSEL 0
`define DP1_11_pad_y 0
`define DP1_12 0
`define DP1_12_GPIO_OUTPUT_ENABLE 0
`define DP1_12_INFUNC_EN 0
`define DP1_12_OUTFUNC_SEL 0
`define DP1_12_PINCTRL_0_IE 0
`define DP1_12_PINCTRL_0_OD 0
`define DP1_12_PULLEN 0
`define DP1_12_PULLSEL 0
`define DP1_12_pad_y 0
`define DP1_13 0
`define DP1_13_GPIO_OUTPUT_ENABLE 0
`define DP1_13_INFUNC_EN 0
`define DP1_13_OUTFUNC_SEL 0
`define DP1_13_PINCTRL_0_IE 0
`define DP1_13_PINCTRL_0_OD 0
`define DP1_13_PULLEN 0
`define DP1_13_PULLSEL 0
`define DP1_13_pad_y 0
`define DP1_14 0
`define DP1_14_GPIO_OUTPUT_ENABLE 0
`define DP1_14_INFUNC_EN 0
`define DP1_14_OUTFUNC_SEL 0
`define DP1_14_PINCTRL_0_IE 0
`define DP1_14_PINCTRL_0_OD 0
`define DP1_14_PULLEN 0
`define DP1_14_PULLSEL 0
`define DP1_14_pad_y 0
`define DP1_15 0
`define DP1_15_GPIO_OUTPUT_ENABLE 0
`define DP1_15_INFUNC_EN 0
`define DP1_15_OUTFUNC_SEL 0
`define DP1_15_PINCTRL_0_IE 0
`define DP1_15_PINCTRL_0_OD 0
`define DP1_15_PULLEN 0
`define DP1_15_PULLSEL 0
`define DP1_15_pad_y 0
`define DP1_16 0
`define DP1_16_GPIO_OUTPUT_ENABLE 0
`define DP1_16_INFUNC_EN 0
`define DP1_16_OUTFUNC_SEL 0
`define DP1_16_PINCTRL_0_IE 0
`define DP1_16_PINCTRL_0_OD 0
`define DP1_16_PULLEN 0
`define DP1_16_PULLSEL 0
`define DP1_16_pad_y 0
`define DP1_17 0
`define DP1_17_GPIO_OUTPUT_ENABLE 0
`define DP1_17_INFUNC_EN 0
`define DP1_17_OUTFUNC_SEL 0
`define DP1_17_PINCTRL_0_IE 0
`define DP1_17_PINCTRL_0_OD 0
`define DP1_17_PULLEN 0
`define DP1_17_PULLSEL 0
`define DP1_17_pad_y 0
`define DP1_18 0
`define DP1_18_GPIO_OUTPUT_ENABLE 0
`define DP1_18_INFUNC_EN 0
`define DP1_18_OUTFUNC_SEL 0
`define DP1_18_PINCTRL_0_IE 0
`define DP1_18_PINCTRL_0_OD 0
`define DP1_18_PULLEN 0
`define DP1_18_PULLSEL 0
`define DP1_18_pad_y 0
`define DP1_19 0
`define DP1_19_GPIO_OUTPUT_ENABLE 0
`define DP1_19_INFUNC_EN 0
`define DP1_19_OUTFUNC_SEL 0
`define DP1_19_PINCTRL_0_IE 0
`define DP1_19_PINCTRL_0_OD 0
`define DP1_19_PULLEN 0
`define DP1_19_PULLSEL 0
`define DP1_19_pad_y 0
`define DP1_1_GPIO_OUTPUT_ENABLE 0
`define DP1_1_INFUNC_EN 0
`define DP1_1_OUTFUNC_SEL 0
`define DP1_1_PINCTRL_0_IE 0
`define DP1_1_PINCTRL_0_OD 0
`define DP1_1_PULLEN 0
`define DP1_1_PULLSEL 0
`define DP1_1_pad_y 0
`define DP1_2 0
`define DP1_20 0
`define DP1_20_GPIO_OUTPUT_ENABLE 0
`define DP1_20_INFUNC_EN 0
`define DP1_20_OUTFUNC_SEL 0
`define DP1_20_PINCTRL_0_IE 0
`define DP1_20_PINCTRL_0_OD 0
`define DP1_20_PULLEN 0
`define DP1_20_PULLSEL 0
`define DP1_20_pad_y 0
`define DP1_21 0
`define DP1_21_GPIO_OUTPUT_ENABLE 0
`define DP1_21_INFUNC_EN 0
`define DP1_21_OUTFUNC_SEL 0
`define DP1_21_PINCTRL_0_IE 0
`define DP1_21_PINCTRL_0_OD 0
`define DP1_21_PULLEN 0
`define DP1_21_PULLSEL 0
`define DP1_21_pad_y 0
`define DP1_22 0
`define DP1_22_GPIO_OUTPUT_ENABLE 0
`define DP1_22_INFUNC_EN 0
`define DP1_22_OUTFUNC_SEL 0
`define DP1_22_PINCTRL_0_IE 0
`define DP1_22_PINCTRL_0_OD 0
`define DP1_22_PULLEN 0
`define DP1_22_PULLSEL 0
`define DP1_22_pad_y 0
`define DP1_23 0
`define DP1_23_GPIO_OUTPUT_ENABLE 0
`define DP1_23_INFUNC_EN 0
`define DP1_23_OUTFUNC_SEL 0
`define DP1_23_PINCTRL_0_IE 0
`define DP1_23_PINCTRL_0_OD 0
`define DP1_23_PULLEN 0
`define DP1_23_PULLSEL 0
`define DP1_23_pad_y 0
`define DP1_24 0
`define DP1_24_GPIO_OUTPUT_ENABLE 0
`define DP1_24_INFUNC_EN 0
`define DP1_24_OUTFUNC_SEL 0
`define DP1_24_PINCTRL_0_IE 0
`define DP1_24_PINCTRL_0_OD 0
`define DP1_24_PULLEN 0
`define DP1_24_PULLSEL 0
`define DP1_24_pad_y 0
`define DP1_25 0
`define DP1_25_GPIO_OUTPUT_ENABLE 0
`define DP1_25_INFUNC_EN 0
`define DP1_25_OUTFUNC_SEL 0
`define DP1_25_PINCTRL_0_IE 0
`define DP1_25_PINCTRL_0_OD 0
`define DP1_25_PULLEN 0
`define DP1_25_PULLSEL 0
`define DP1_25_pad_y 0
`define DP1_26 0
`define DP1_26_GPIO_OUTPUT_ENABLE 0
`define DP1_26_INFUNC_EN 0
`define DP1_26_OUTFUNC_SEL 0
`define DP1_26_PINCTRL_0_IE 0
`define DP1_26_PINCTRL_0_OD 0
`define DP1_26_PULLEN 0
`define DP1_26_PULLSEL 0
`define DP1_26_pad_y 0
`define DP1_27 0
`define DP1_27_GPIO_OUTPUT_ENABLE 0
`define DP1_27_INFUNC_EN 0
`define DP1_27_OUTFUNC_SEL 0
`define DP1_27_PINCTRL_0_IE 0
`define DP1_27_PINCTRL_0_OD 0
`define DP1_27_PULLEN 0
`define DP1_27_PULLSEL 0
`define DP1_27_pad_y 0
`define DP1_28 0
`define DP1_28_GPIO_OUTPUT_ENABLE 0
`define DP1_28_INFUNC_EN 0
`define DP1_28_OUTFUNC_SEL 0
`define DP1_28_PINCTRL_0_IE 0
`define DP1_28_PINCTRL_0_OD 0
`define DP1_28_PULLEN 0
`define DP1_28_PULLSEL 0
`define DP1_28_pad_y 0
`define DP1_29 0
`define DP1_29_GPIO_OUTPUT_ENABLE 0
`define DP1_29_INFUNC_EN 0
`define DP1_29_OUTFUNC_SEL 0
`define DP1_29_PINCTRL_0_IE 0
`define DP1_29_PINCTRL_0_OD 0
`define DP1_29_PULLEN 0
`define DP1_29_PULLSEL 0
`define DP1_29_pad_y 0
`define DP1_2_GPIO_OUTPUT_ENABLE 0
`define DP1_2_INFUNC_EN 0
`define DP1_2_OUTFUNC_SEL 0
`define DP1_2_PINCTRL_0_IE 0
`define DP1_2_PINCTRL_0_OD 0
`define DP1_2_PULLEN 0
`define DP1_2_PULLSEL 0
`define DP1_2_pad_y 0
`define DP1_3 0
`define DP1_30 0
`define DP1_30_GPIO_OUTPUT_ENABLE 0
`define DP1_30_INFUNC_EN 0
`define DP1_30_OUTFUNC_SEL 0
`define DP1_30_PINCTRL_0_IE 0
`define DP1_30_PINCTRL_0_OD 0
`define DP1_30_PULLEN 0
`define DP1_30_PULLSEL 0
`define DP1_30_pad_y 0
`define DP1_31 0
`define DP1_31_GPIO_OUTPUT_ENABLE 0
`define DP1_31_INFUNC_EN 0
`define DP1_31_OUTFUNC_SEL 0
`define DP1_31_PINCTRL_0_IE 0
`define DP1_31_PINCTRL_0_OD 0
`define DP1_31_PULLEN 0
`define DP1_31_PULLSEL 0
`define DP1_31_pad_y 0
`define DP1_3_GPIO_OUTPUT_ENABLE 0
`define DP1_3_INFUNC_EN 0
`define DP1_3_OUTFUNC_SEL 0
`define DP1_3_PINCTRL_0_IE 0
`define DP1_3_PINCTRL_0_OD 0
`define DP1_3_PULLEN 0
`define DP1_3_PULLSEL 0
`define DP1_3_pad_y 0
`define DP1_4 0
`define DP1_4_GPIO_OUTPUT_ENABLE 0
`define DP1_4_INFUNC_EN 0
`define DP1_4_OUTFUNC_SEL 0
`define DP1_4_PINCTRL_0_IE 0
`define DP1_4_PINCTRL_0_OD 0
`define DP1_4_PULLEN 0
`define DP1_4_PULLSEL 0
`define DP1_4_pad_y 0
`define DP1_5 0
`define DP1_5_GPIO_OUTPUT_ENABLE 0
`define DP1_5_INFUNC_EN 0
`define DP1_5_OUTFUNC_SEL 0
`define DP1_5_PINCTRL_0_IE 0
`define DP1_5_PINCTRL_0_OD 0
`define DP1_5_PULLEN 0
`define DP1_5_PULLSEL 0
`define DP1_5_pad_y 0
`define DP1_6 0
`define DP1_6_GPIO_OUTPUT_ENABLE 0
`define DP1_6_INFUNC_EN 0
`define DP1_6_OUTFUNC_SEL 0
`define DP1_6_PINCTRL_0_IE 0
`define DP1_6_PINCTRL_0_OD 0
`define DP1_6_PULLEN 0
`define DP1_6_PULLSEL 0
`define DP1_6_pad_y 0
`define DP1_7 0
`define DP1_7_GPIO_OUTPUT_ENABLE 0
`define DP1_7_INFUNC_EN 0
`define DP1_7_OUTFUNC_SEL 0
`define DP1_7_PINCTRL_0_IE 0
`define DP1_7_PINCTRL_0_OD 0
`define DP1_7_PULLEN 0
`define DP1_7_PULLSEL 0
`define DP1_7_pad_y 0
`define DP1_8 0
`define DP1_8_GPIO_OUTPUT_ENABLE 0
`define DP1_8_INFUNC_EN 0
`define DP1_8_OUTFUNC_SEL 0
`define DP1_8_PINCTRL_0_IE 0
`define DP1_8_PINCTRL_0_OD 0
`define DP1_8_PULLEN 0
`define DP1_8_PULLSEL 0
`define DP1_8_pad_y 0
`define DP1_9 0
`define DP1_9_GPIO_OUTPUT_ENABLE 0
`define DP1_9_INFUNC_EN 0
`define DP1_9_OUTFUNC_SEL 0
`define DP1_9_PINCTRL_0_IE 0
`define DP1_9_PINCTRL_0_OD 0
`define DP1_9_PULLEN 0
`define DP1_9_PULLSEL 0
`define DP1_9_pad_y 0
`define DP2_0 0
`define DP2_0_GPIO_OUTPUT_ENABLE 0
`define DP2_0_INFUNC_EN 0
`define DP2_0_OUTFUNC_SEL 0
`define DP2_0_PINCTRL_0_IE 0
`define DP2_0_PINCTRL_0_OD 0
`define DP2_0_PULLEN 0
`define DP2_0_PULLSEL 0
`define DP2_0_pad_y 0
`define DP2_1 0
`define DP2_10 0
`define DP2_10_GPIO_OUTPUT_ENABLE 0
`define DP2_10_INFUNC_EN 0
`define DP2_10_OUTFUNC_SEL 0
`define DP2_10_PINCTRL_0_IE 0
`define DP2_10_PINCTRL_0_OD 0
`define DP2_10_PULLEN 0
`define DP2_10_PULLSEL 0
`define DP2_10_pad_y 0
`define DP2_11 0
`define DP2_11_GPIO_OUTPUT_ENABLE 0
`define DP2_11_INFUNC_EN 0
`define DP2_11_OUTFUNC_SEL 0
`define DP2_11_PINCTRL_0_IE 0
`define DP2_11_PINCTRL_0_OD 0
`define DP2_11_PULLEN 0
`define DP2_11_PULLSEL 0
`define DP2_11_pad_y 0
`define DP2_12 0
`define DP2_12_GPIO_OUTPUT_ENABLE 0
`define DP2_12_INFUNC_EN 0
`define DP2_12_OUTFUNC_SEL 0
`define DP2_12_PINCTRL_0_IE 0
`define DP2_12_PINCTRL_0_OD 0
`define DP2_12_PULLEN 0
`define DP2_12_PULLSEL 0
`define DP2_12_pad_y 0
`define DP2_13 0
`define DP2_13_GPIO_OUTPUT_ENABLE 0
`define DP2_13_INFUNC_EN 0
`define DP2_13_OUTFUNC_SEL 0
`define DP2_13_PINCTRL_0_IE 0
`define DP2_13_PINCTRL_0_OD 0
`define DP2_13_PULLEN 0
`define DP2_13_PULLSEL 0
`define DP2_13_pad_y 0
`define DP2_14 0
`define DP2_14_GPIO_OUTPUT_ENABLE 0
`define DP2_14_INFUNC_EN 0
`define DP2_14_OUTFUNC_SEL 0
`define DP2_14_PINCTRL_0_IE 0
`define DP2_14_PINCTRL_0_OD 0
`define DP2_14_PULLEN 0
`define DP2_14_PULLSEL 0
`define DP2_14_pad_y 0
`define DP2_15 0
`define DP2_15_GPIO_OUTPUT_ENABLE 0
`define DP2_15_INFUNC_EN 0
`define DP2_15_OUTFUNC_SEL 0
`define DP2_15_PINCTRL_0_IE 0
`define DP2_15_PINCTRL_0_OD 0
`define DP2_15_PULLEN 0
`define DP2_15_PULLSEL 0
`define DP2_15_pad_y 0
`define DP2_16 0
`define DP2_16_GPIO_OUTPUT_ENABLE 0
`define DP2_16_INFUNC_EN 0
`define DP2_16_OUTFUNC_SEL 0
`define DP2_16_PINCTRL_0_IE 0
`define DP2_16_PINCTRL_0_OD 0
`define DP2_16_PULLEN 0
`define DP2_16_PULLSEL 0
`define DP2_16_pad_y 0
`define DP2_17 0
`define DP2_17_GPIO_OUTPUT_ENABLE 0
`define DP2_17_INFUNC_EN 0
`define DP2_17_OUTFUNC_SEL 0
`define DP2_17_PINCTRL_0_IE 0
`define DP2_17_PINCTRL_0_OD 0
`define DP2_17_PULLEN 0
`define DP2_17_PULLSEL 0
`define DP2_17_pad_y 0
`define DP2_18 0
`define DP2_18_GPIO_OUTPUT_ENABLE 0
`define DP2_18_INFUNC_EN 0
`define DP2_18_OUTFUNC_SEL 0
`define DP2_18_PINCTRL_0_IE 0
`define DP2_18_PINCTRL_0_OD 0
`define DP2_18_PULLEN 0
`define DP2_18_PULLSEL 0
`define DP2_18_pad_y 0
`define DP2_19 0
`define DP2_19_GPIO_OUTPUT_ENABLE 0
`define DP2_19_INFUNC_EN 0
`define DP2_19_OUTFUNC_SEL 0
`define DP2_19_PINCTRL_0_IE 0
`define DP2_19_PINCTRL_0_OD 0
`define DP2_19_PULLEN 0
`define DP2_19_PULLSEL 0
`define DP2_19_pad_y 0
`define DP2_1_GPIO_OUTPUT_ENABLE 0
`define DP2_1_INFUNC_EN 0
`define DP2_1_OUTFUNC_SEL 0
`define DP2_1_PINCTRL_0_IE 0
`define DP2_1_PINCTRL_0_OD 0
`define DP2_1_PULLEN 0
`define DP2_1_PULLSEL 0
`define DP2_1_pad_y 0
`define DP2_2 0
`define DP2_20 0
`define DP2_20_GPIO_OUTPUT_ENABLE 0
`define DP2_20_INFUNC_EN 0
`define DP2_20_OUTFUNC_SEL 0
`define DP2_20_PINCTRL_0_IE 0
`define DP2_20_PINCTRL_0_OD 0
`define DP2_20_PULLEN 0
`define DP2_20_PULLSEL 0
`define DP2_20_pad_y 0
`define DP2_21 0
`define DP2_21_GPIO_OUTPUT_ENABLE 0
`define DP2_21_INFUNC_EN 0
`define DP2_21_OUTFUNC_SEL 0
`define DP2_21_PINCTRL_0_IE 0
`define DP2_21_PINCTRL_0_OD 0
`define DP2_21_PULLEN 0
`define DP2_21_PULLSEL 0
`define DP2_21_pad_y 0
`define DP2_22 0
`define DP2_22_GPIO_OUTPUT_ENABLE 0
`define DP2_22_INFUNC_EN 0
`define DP2_22_OUTFUNC_SEL 0
`define DP2_22_PINCTRL_0_IE 0
`define DP2_22_PINCTRL_0_OD 0
`define DP2_22_PULLEN 0
`define DP2_22_PULLSEL 0
`define DP2_22_pad_y 0
`define DP2_23 0
`define DP2_23_GPIO_OUTPUT_ENABLE 0
`define DP2_23_INFUNC_EN 0
`define DP2_23_OUTFUNC_SEL 0
`define DP2_23_PINCTRL_0_IE 0
`define DP2_23_PINCTRL_0_OD 0
`define DP2_23_PULLEN 0
`define DP2_23_PULLSEL 0
`define DP2_23_pad_y 0
`define DP2_24 0
`define DP2_24_GPIO_OUTPUT_ENABLE 0
`define DP2_24_INFUNC_EN 0
`define DP2_24_OUTFUNC_SEL 0
`define DP2_24_PINCTRL_0_IE 0
`define DP2_24_PINCTRL_0_OD 0
`define DP2_24_PULLEN 0
`define DP2_24_PULLSEL 0
`define DP2_24_pad_y 0
`define DP2_25 0
`define DP2_25_GPIO_OUTPUT_ENABLE 0
`define DP2_25_INFUNC_EN 0
`define DP2_25_OUTFUNC_SEL 0
`define DP2_25_PINCTRL_0_IE 0
`define DP2_25_PINCTRL_0_OD 0
`define DP2_25_PULLEN 0
`define DP2_25_PULLSEL 0
`define DP2_25_pad_y 0
`define DP2_26 0
`define DP2_26_GPIO_OUTPUT_ENABLE 0
`define DP2_26_INFUNC_EN 0
`define DP2_26_OUTFUNC_SEL 0
`define DP2_26_PINCTRL_0_IE 0
`define DP2_26_PINCTRL_0_OD 0
`define DP2_26_PULLEN 0
`define DP2_26_PULLSEL 0
`define DP2_26_pad_y 0
`define DP2_27 0
`define DP2_27_GPIO_OUTPUT_ENABLE 0
`define DP2_27_INFUNC_EN 0
`define DP2_27_OUTFUNC_SEL 0
`define DP2_27_PINCTRL_0_IE 0
`define DP2_27_PINCTRL_0_OD 0
`define DP2_27_PULLEN 0
`define DP2_27_PULLSEL 0
`define DP2_27_pad_y 0
`define DP2_28 0
`define DP2_28_GPIO_OUTPUT_ENABLE 0
`define DP2_28_INFUNC_EN 0
`define DP2_28_OUTFUNC_SEL 0
`define DP2_28_PINCTRL_0_IE 0
`define DP2_28_PINCTRL_0_OD 0
`define DP2_28_PULLEN 0
`define DP2_28_PULLSEL 0
`define DP2_28_pad_y 0
`define DP2_29 0
`define DP2_29_GPIO_OUTPUT_ENABLE 0
`define DP2_29_INFUNC_EN 0
`define DP2_29_OUTFUNC_SEL 0
`define DP2_29_PINCTRL_0_IE 0
`define DP2_29_PINCTRL_0_OD 0
`define DP2_29_PULLEN 0
`define DP2_29_PULLSEL 0
`define DP2_29_pad_y 0
`define DP2_2_GPIO_OUTPUT_ENABLE 0
`define DP2_2_INFUNC_EN 0
`define DP2_2_OUTFUNC_SEL 0
`define DP2_2_PINCTRL_0_IE 0
`define DP2_2_PINCTRL_0_OD 0
`define DP2_2_PULLEN 0
`define DP2_2_PULLSEL 0
`define DP2_2_pad_y 0
`define DP2_3 0
`define DP2_30 0
`define DP2_30_GPIO_OUTPUT_ENABLE 0
`define DP2_30_INFUNC_EN 0
`define DP2_30_OUTFUNC_SEL 0
`define DP2_30_PINCTRL_0_IE 0
`define DP2_30_PINCTRL_0_OD 0
`define DP2_30_PULLEN 0
`define DP2_30_PULLSEL 0
`define DP2_30_pad_y 0
`define DP2_31 0
`define DP2_31_GPIO_OUTPUT_ENABLE 0
`define DP2_31_INFUNC_EN 0
`define DP2_31_OUTFUNC_SEL 0
`define DP2_31_PINCTRL_0_IE 0
`define DP2_31_PINCTRL_0_OD 0
`define DP2_31_PULLEN 0
`define DP2_31_PULLSEL 0
`define DP2_31_pad_y 0
`define DP2_3_GPIO_OUTPUT_ENABLE 0
`define DP2_3_INFUNC_EN 0
`define DP2_3_OUTFUNC_SEL 0
`define DP2_3_PINCTRL_0_IE 0
`define DP2_3_PINCTRL_0_OD 0
`define DP2_3_PULLEN 0
`define DP2_3_PULLSEL 0
`define DP2_3_pad_y 0
`define DP2_4 0
`define DP2_4_GPIO_OUTPUT_ENABLE 0
`define DP2_4_INFUNC_EN 0
`define DP2_4_OUTFUNC_SEL 0
`define DP2_4_PINCTRL_0_IE 0
`define DP2_4_PINCTRL_0_OD 0
`define DP2_4_PULLEN 0
`define DP2_4_PULLSEL 0
`define DP2_4_pad_y 0
`define DP2_5 0
`define DP2_5_GPIO_OUTPUT_ENABLE 0
`define DP2_5_INFUNC_EN 0
`define DP2_5_OUTFUNC_SEL 0
`define DP2_5_PINCTRL_0_IE 0
`define DP2_5_PINCTRL_0_OD 0
`define DP2_5_PULLEN 0
`define DP2_5_PULLSEL 0
`define DP2_5_pad_y 0
`define DP2_6 0
`define DP2_6_GPIO_OUTPUT_ENABLE 0
`define DP2_6_INFUNC_EN 0
`define DP2_6_OUTFUNC_SEL 0
`define DP2_6_PINCTRL_0_IE 0
`define DP2_6_PINCTRL_0_OD 0
`define DP2_6_PULLEN 0
`define DP2_6_PULLSEL 0
`define DP2_6_pad_y 0
`define DP2_7 0
`define DP2_7_GPIO_OUTPUT_ENABLE 0
`define DP2_7_INFUNC_EN 0
`define DP2_7_OUTFUNC_SEL 0
`define DP2_7_PINCTRL_0_IE 0
`define DP2_7_PINCTRL_0_OD 0
`define DP2_7_PULLEN 0
`define DP2_7_PULLSEL 0
`define DP2_7_pad_y 0
`define DP2_8 0
`define DP2_8_GPIO_OUTPUT_ENABLE 0
`define DP2_8_INFUNC_EN 0
`define DP2_8_OUTFUNC_SEL 0
`define DP2_8_PINCTRL_0_IE 0
`define DP2_8_PINCTRL_0_OD 0
`define DP2_8_PULLEN 0
`define DP2_8_PULLSEL 0
`define DP2_8_pad_y 0
`define DP2_9 0
`define DP2_9_GPIO_OUTPUT_ENABLE 0
`define DP2_9_INFUNC_EN 0
`define DP2_9_OUTFUNC_SEL 0
`define DP2_9_PINCTRL_0_IE 0
`define DP2_9_PINCTRL_0_OD 0
`define DP2_9_PULLEN 0
`define DP2_9_PULLSEL 0
`define DP2_9_pad_y 0
`define DP3_0 0
`define DP3_0_GPIO_OUTPUT_ENABLE 0
`define DP3_0_INFUNC_EN 0
`define DP3_0_OUTFUNC_SEL 0
`define DP3_0_PINCTRL_0_IE 0
`define DP3_0_PINCTRL_0_OD 0
`define DP3_0_PULLEN 0
`define DP3_0_PULLSEL 0
`define DP3_0_pad_y 0
`define DP3_1 0
`define DP3_10 0
`define DP3_10_GPIO_OUTPUT_ENABLE 0
`define DP3_10_INFUNC_EN 0
`define DP3_10_OUTFUNC_SEL 0
`define DP3_10_PINCTRL_0_IE 0
`define DP3_10_PINCTRL_0_OD 0
`define DP3_10_PULLEN 0
`define DP3_10_PULLSEL 0
`define DP3_10_pad_y 0
`define DP3_11 0
`define DP3_11_GPIO_OUTPUT_ENABLE 0
`define DP3_11_INFUNC_EN 0
`define DP3_11_OUTFUNC_SEL 0
`define DP3_11_PINCTRL_0_IE 0
`define DP3_11_PINCTRL_0_OD 0
`define DP3_11_PULLEN 0
`define DP3_11_PULLSEL 0
`define DP3_11_pad_y 0
`define DP3_12 0
`define DP3_12_GPIO_OUTPUT_ENABLE 0
`define DP3_12_INFUNC_EN 0
`define DP3_12_OUTFUNC_SEL 0
`define DP3_12_PINCTRL_0_IE 0
`define DP3_12_PINCTRL_0_OD 0
`define DP3_12_PULLEN 0
`define DP3_12_PULLSEL 0
`define DP3_12_pad_y 0
`define DP3_13 0
`define DP3_13_GPIO_OUTPUT_ENABLE 0
`define DP3_13_INFUNC_EN 0
`define DP3_13_OUTFUNC_SEL 0
`define DP3_13_PINCTRL_0_IE 0
`define DP3_13_PINCTRL_0_OD 0
`define DP3_13_PULLEN 0
`define DP3_13_PULLSEL 0
`define DP3_13_pad_y 0
`define DP3_14 0
`define DP3_14_GPIO_OUTPUT_ENABLE 0
`define DP3_14_INFUNC_EN 0
`define DP3_14_OUTFUNC_SEL 0
`define DP3_14_PINCTRL_0_IE 0
`define DP3_14_PINCTRL_0_OD 0
`define DP3_14_PULLEN 0
`define DP3_14_PULLSEL 0
`define DP3_14_pad_y 0
`define DP3_15 0
`define DP3_15_GPIO_OUTPUT_ENABLE 0
`define DP3_15_INFUNC_EN 0
`define DP3_15_OUTFUNC_SEL 0
`define DP3_15_PINCTRL_0_IE 0
`define DP3_15_PINCTRL_0_OD 0
`define DP3_15_PULLEN 0
`define DP3_15_PULLSEL 0
`define DP3_15_pad_y 0
`define DP3_16 0
`define DP3_16_GPIO_OUTPUT_ENABLE 0
`define DP3_16_INFUNC_EN 0
`define DP3_16_OUTFUNC_SEL 0
`define DP3_16_PINCTRL_0_IE 0
`define DP3_16_PINCTRL_0_OD 0
`define DP3_16_PULLEN 0
`define DP3_16_PULLSEL 0
`define DP3_16_pad_y 0
`define DP3_17 0
`define DP3_17_GPIO_OUTPUT_ENABLE 0
`define DP3_17_INFUNC_EN 0
`define DP3_17_OUTFUNC_SEL 0
`define DP3_17_PINCTRL_0_IE 0
`define DP3_17_PINCTRL_0_OD 0
`define DP3_17_PULLEN 0
`define DP3_17_PULLSEL 0
`define DP3_17_pad_y 0
`define DP3_18 0
`define DP3_18_GPIO_OUTPUT_ENABLE 0
`define DP3_18_INFUNC_EN 0
`define DP3_18_OUTFUNC_SEL 0
`define DP3_18_PINCTRL_0_IE 0
`define DP3_18_PINCTRL_0_OD 0
`define DP3_18_PULLEN 0
`define DP3_18_PULLSEL 0
`define DP3_18_pad_y 0
`define DP3_19 0
`define DP3_19_GPIO_OUTPUT_ENABLE 0
`define DP3_19_INFUNC_EN 0
`define DP3_19_OUTFUNC_SEL 0
`define DP3_19_PINCTRL_0_IE 0
`define DP3_19_PINCTRL_0_OD 0
`define DP3_19_PULLEN 0
`define DP3_19_PULLSEL 0
`define DP3_19_pad_y 0
`define DP3_1_GPIO_OUTPUT_ENABLE 0
`define DP3_1_INFUNC_EN 0
`define DP3_1_OUTFUNC_SEL 0
`define DP3_1_PINCTRL_0_IE 0
`define DP3_1_PINCTRL_0_OD 0
`define DP3_1_PULLEN 0
`define DP3_1_PULLSEL 0
`define DP3_1_pad_y 0
`define DP3_2 0
`define DP3_20 0
`define DP3_20_GPIO_OUTPUT_ENABLE 0
`define DP3_20_INFUNC_EN 0
`define DP3_20_OUTFUNC_SEL 0
`define DP3_20_PINCTRL_0_IE 0
`define DP3_20_PINCTRL_0_OD 0
`define DP3_20_PULLEN 0
`define DP3_20_PULLSEL 0
`define DP3_20_pad_y 0
`define DP3_21 0
`define DP3_21_GPIO_OUTPUT_ENABLE 0
`define DP3_21_INFUNC_EN 0
`define DP3_21_OUTFUNC_SEL 0
`define DP3_21_PINCTRL_0_IE 0
`define DP3_21_PINCTRL_0_OD 0
`define DP3_21_PULLEN 0
`define DP3_21_PULLSEL 0
`define DP3_21_pad_y 0
`define DP3_22 0
`define DP3_22_GPIO_OUTPUT_ENABLE 0
`define DP3_22_INFUNC_EN 0
`define DP3_22_OUTFUNC_SEL 0
`define DP3_22_PINCTRL_0_IE 0
`define DP3_22_PINCTRL_0_OD 0
`define DP3_22_PULLEN 0
`define DP3_22_PULLSEL 0
`define DP3_22_pad_y 0
`define DP3_23 0
`define DP3_23_GPIO_OUTPUT_ENABLE 0
`define DP3_23_INFUNC_EN 0
`define DP3_23_OUTFUNC_SEL 0
`define DP3_23_PINCTRL_0_IE 0
`define DP3_23_PINCTRL_0_OD 0
`define DP3_23_PULLEN 0
`define DP3_23_PULLSEL 0
`define DP3_23_pad_y 0
`define DP3_24 0
`define DP3_24_GPIO_OUTPUT_ENABLE 0
`define DP3_24_INFUNC_EN 0
`define DP3_24_OUTFUNC_SEL 0
`define DP3_24_PINCTRL_0_IE 0
`define DP3_24_PINCTRL_0_OD 0
`define DP3_24_PULLEN 0
`define DP3_24_PULLSEL 0
`define DP3_24_pad_y 0
`define DP3_25 0
`define DP3_25_GPIO_OUTPUT_ENABLE 0
`define DP3_25_INFUNC_EN 0
`define DP3_25_OUTFUNC_SEL 0
`define DP3_25_PINCTRL_0_IE 0
`define DP3_25_PINCTRL_0_OD 0
`define DP3_25_PULLEN 0
`define DP3_25_PULLSEL 0
`define DP3_25_pad_y 0
`define DP3_26 0
`define DP3_26_GPIO_OUTPUT_ENABLE 0
`define DP3_26_INFUNC_EN 0
`define DP3_26_OUTFUNC_SEL 0
`define DP3_26_PINCTRL_0_IE 0
`define DP3_26_PINCTRL_0_OD 0
`define DP3_26_PULLEN 0
`define DP3_26_PULLSEL 0
`define DP3_26_pad_y 0
`define DP3_27 0
`define DP3_27_GPIO_OUTPUT_ENABLE 0
`define DP3_27_INFUNC_EN 0
`define DP3_27_OUTFUNC_SEL 0
`define DP3_27_PINCTRL_0_IE 0
`define DP3_27_PINCTRL_0_OD 0
`define DP3_27_PULLEN 0
`define DP3_27_PULLSEL 0
`define DP3_27_pad_y 0
`define DP3_28 0
`define DP3_28_GPIO_OUTPUT_ENABLE 0
`define DP3_28_INFUNC_EN 0
`define DP3_28_OUTFUNC_SEL 0
`define DP3_28_PINCTRL_0_IE 0
`define DP3_28_PINCTRL_0_OD 0
`define DP3_28_PULLEN 0
`define DP3_28_PULLSEL 0
`define DP3_28_pad_y 0
`define DP3_29 0
`define DP3_29_GPIO_OUTPUT_ENABLE 0
`define DP3_29_INFUNC_EN 0
`define DP3_29_OUTFUNC_SEL 0
`define DP3_29_PINCTRL_0_IE 0
`define DP3_29_PINCTRL_0_OD 0
`define DP3_29_PULLEN 0
`define DP3_29_PULLSEL 0
`define DP3_29_pad_y 0
`define DP3_2_GPIO_OUTPUT_ENABLE 0
`define DP3_2_INFUNC_EN 0
`define DP3_2_OUTFUNC_SEL 0
`define DP3_2_PINCTRL_0_IE 0
`define DP3_2_PINCTRL_0_OD 0
`define DP3_2_PULLEN 0
`define DP3_2_PULLSEL 0
`define DP3_2_pad_y 0
`define DP3_3 0
`define DP3_30 0
`define DP3_30_GPIO_OUTPUT_ENABLE 0
`define DP3_30_INFUNC_EN 0
`define DP3_30_OUTFUNC_SEL 0
`define DP3_30_PINCTRL_0_IE 0
`define DP3_30_PINCTRL_0_OD 0
`define DP3_30_PULLEN 0
`define DP3_30_PULLSEL 0
`define DP3_30_pad_y 0
`define DP3_31 0
`define DP3_31_GPIO_OUTPUT_ENABLE 0
`define DP3_31_INFUNC_EN 0
`define DP3_31_OUTFUNC_SEL 0
`define DP3_31_PINCTRL_0_IE 0
`define DP3_31_PINCTRL_0_OD 0
`define DP3_31_PULLEN 0
`define DP3_31_PULLSEL 0
`define DP3_31_pad_y 0
`define DP3_3_GPIO_OUTPUT_ENABLE 0
`define DP3_3_INFUNC_EN 0
`define DP3_3_OUTFUNC_SEL 0
`define DP3_3_PINCTRL_0_IE 0
`define DP3_3_PINCTRL_0_OD 0
`define DP3_3_PULLEN 0
`define DP3_3_PULLSEL 0
`define DP3_3_pad_y 0
`define DP3_4 0
`define DP3_4_GPIO_OUTPUT_ENABLE 0
`define DP3_4_INFUNC_EN 0
`define DP3_4_OUTFUNC_SEL 0
`define DP3_4_PINCTRL_0_IE 0
`define DP3_4_PINCTRL_0_OD 0
`define DP3_4_PULLEN 0
`define DP3_4_PULLSEL 0
`define DP3_4_pad_y 0
`define DP3_5 0
`define DP3_5_GPIO_OUTPUT_ENABLE 0
`define DP3_5_INFUNC_EN 0
`define DP3_5_OUTFUNC_SEL 0
`define DP3_5_PINCTRL_0_IE 0
`define DP3_5_PINCTRL_0_OD 0
`define DP3_5_PULLEN 0
`define DP3_5_PULLSEL 0
`define DP3_5_pad_y 0
`define DP3_6 0
`define DP3_6_GPIO_OUTPUT_ENABLE 0
`define DP3_6_INFUNC_EN 0
`define DP3_6_OUTFUNC_SEL 0
`define DP3_6_PINCTRL_0_IE 0
`define DP3_6_PINCTRL_0_OD 0
`define DP3_6_PULLEN 0
`define DP3_6_PULLSEL 0
`define DP3_6_pad_y 0
`define DP3_7 0
`define DP3_7_GPIO_OUTPUT_ENABLE 0
`define DP3_7_INFUNC_EN 0
`define DP3_7_OUTFUNC_SEL 0
`define DP3_7_PINCTRL_0_IE 0
`define DP3_7_PINCTRL_0_OD 0
`define DP3_7_PULLEN 0
`define DP3_7_PULLSEL 0
`define DP3_7_pad_y 0
`define DP3_8 0
`define DP3_8_GPIO_OUTPUT_ENABLE 0
`define DP3_8_INFUNC_EN 0
`define DP3_8_OUTFUNC_SEL 0
`define DP3_8_PINCTRL_0_IE 0
`define DP3_8_PINCTRL_0_OD 0
`define DP3_8_PULLEN 0
`define DP3_8_PULLSEL 0
`define DP3_8_pad_y 0
`define DP3_9 0
`define DP3_9_GPIO_OUTPUT_ENABLE 0
`define DP3_9_INFUNC_EN 0
`define DP3_9_OUTFUNC_SEL 0
`define DP3_9_PINCTRL_0_IE 0
`define DP3_9_PINCTRL_0_OD 0
`define DP3_9_PULLEN 0
`define DP3_9_PULLSEL 0
`define DP3_9_pad_y 0
`define DP4_0 0
`define DP4_0_GPIO_OUTPUT_ENABLE 0
`define DP4_0_INFUNC_EN 0
`define DP4_0_OUTFUNC_SEL 0
`define DP4_0_PINCTRL_0_IE 0
`define DP4_0_PINCTRL_0_OD 0
`define DP4_0_PULLEN 0
`define DP4_0_PULLSEL 0
`define DP4_0_pad_y 0
`define DP4_1 0
`define DP4_10 0
`define DP4_10_GPIO_OUTPUT_ENABLE 0
`define DP4_10_INFUNC_EN 0
`define DP4_10_OUTFUNC_SEL 0
`define DP4_10_PINCTRL_0_IE 0
`define DP4_10_PINCTRL_0_OD 0
`define DP4_10_PULLEN 0
`define DP4_10_PULLSEL 0
`define DP4_10_pad_y 0
`define DP4_11 0
`define DP4_11_GPIO_OUTPUT_ENABLE 0
`define DP4_11_INFUNC_EN 0
`define DP4_11_OUTFUNC_SEL 0
`define DP4_11_PINCTRL_0_IE 0
`define DP4_11_PINCTRL_0_OD 0
`define DP4_11_PULLEN 0
`define DP4_11_PULLSEL 0
`define DP4_11_pad_y 0
`define DP4_12 0
`define DP4_12_GPIO_OUTPUT_ENABLE 0
`define DP4_12_INFUNC_EN 0
`define DP4_12_OUTFUNC_SEL 0
`define DP4_12_PINCTRL_0_IE 0
`define DP4_12_PINCTRL_0_OD 0
`define DP4_12_PULLEN 0
`define DP4_12_PULLSEL 0
`define DP4_12_pad_y 0
`define DP4_13 0
`define DP4_13_GPIO_OUTPUT_ENABLE 0
`define DP4_13_INFUNC_EN 0
`define DP4_13_OUTFUNC_SEL 0
`define DP4_13_PINCTRL_0_IE 0
`define DP4_13_PINCTRL_0_OD 0
`define DP4_13_PULLEN 0
`define DP4_13_PULLSEL 0
`define DP4_13_pad_y 0
`define DP4_14 0
`define DP4_14_GPIO_OUTPUT_ENABLE 0
`define DP4_14_INFUNC_EN 0
`define DP4_14_OUTFUNC_SEL 0
`define DP4_14_PINCTRL_0_IE 0
`define DP4_14_PINCTRL_0_OD 0
`define DP4_14_PULLEN 0
`define DP4_14_PULLSEL 0
`define DP4_14_pad_y 0
`define DP4_15 0
`define DP4_15_GPIO_OUTPUT_ENABLE 0
`define DP4_15_INFUNC_EN 0
`define DP4_15_OUTFUNC_SEL 0
`define DP4_15_PINCTRL_0_IE 0
`define DP4_15_PINCTRL_0_OD 0
`define DP4_15_PULLEN 0
`define DP4_15_PULLSEL 0
`define DP4_15_pad_y 0
`define DP4_16 0
`define DP4_16_GPIO_OUTPUT_ENABLE 0
`define DP4_16_INFUNC_EN 0
`define DP4_16_OUTFUNC_SEL 0
`define DP4_16_PINCTRL_0_IE 0
`define DP4_16_PINCTRL_0_OD 0
`define DP4_16_PULLEN 0
`define DP4_16_PULLSEL 0
`define DP4_16_pad_y 0
`define DP4_17 0
`define DP4_17_GPIO_OUTPUT_ENABLE 0
`define DP4_17_INFUNC_EN 0
`define DP4_17_OUTFUNC_SEL 0
`define DP4_17_PINCTRL_0_IE 0
`define DP4_17_PINCTRL_0_OD 0
`define DP4_17_PULLEN 0
`define DP4_17_PULLSEL 0
`define DP4_17_pad_y 0
`define DP4_18 0
`define DP4_18_GPIO_OUTPUT_ENABLE 0
`define DP4_18_INFUNC_EN 0
`define DP4_18_OUTFUNC_SEL 0
`define DP4_18_PINCTRL_0_IE 0
`define DP4_18_PINCTRL_0_OD 0
`define DP4_18_PULLEN 0
`define DP4_18_PULLSEL 0
`define DP4_18_pad_y 0
`define DP4_19 0
`define DP4_19_GPIO_OUTPUT_ENABLE 0
`define DP4_19_INFUNC_EN 0
`define DP4_19_OUTFUNC_SEL 0
`define DP4_19_PINCTRL_0_IE 0
`define DP4_19_PINCTRL_0_OD 0
`define DP4_19_PULLEN 0
`define DP4_19_PULLSEL 0
`define DP4_19_pad_y 0
`define DP4_1_GPIO_OUTPUT_ENABLE 0
`define DP4_1_INFUNC_EN 0
`define DP4_1_OUTFUNC_SEL 0
`define DP4_1_PINCTRL_0_IE 0
`define DP4_1_PINCTRL_0_OD 0
`define DP4_1_PULLEN 0
`define DP4_1_PULLSEL 0
`define DP4_1_pad_y 0
`define DP4_2 0
`define DP4_20 0
`define DP4_20_GPIO_OUTPUT_ENABLE 0
`define DP4_20_INFUNC_EN 0
`define DP4_20_OUTFUNC_SEL 0
`define DP4_20_PINCTRL_0_IE 0
`define DP4_20_PINCTRL_0_OD 0
`define DP4_20_PULLEN 0
`define DP4_20_PULLSEL 0
`define DP4_20_pad_y 0
`define DP4_21 0
`define DP4_21_GPIO_OUTPUT_ENABLE 0
`define DP4_21_INFUNC_EN 0
`define DP4_21_OUTFUNC_SEL 0
`define DP4_21_PINCTRL_0_IE 0
`define DP4_21_PINCTRL_0_OD 0
`define DP4_21_PULLEN 0
`define DP4_21_PULLSEL 0
`define DP4_21_pad_y 0
`define DP4_22 0
`define DP4_22_GPIO_OUTPUT_ENABLE 0
`define DP4_22_INFUNC_EN 0
`define DP4_22_OUTFUNC_SEL 0
`define DP4_22_PINCTRL_0_IE 0
`define DP4_22_PINCTRL_0_OD 0
`define DP4_22_PULLEN 0
`define DP4_22_PULLSEL 0
`define DP4_22_pad_y 0
`define DP4_23 0
`define DP4_23_GPIO_OUTPUT_ENABLE 0
`define DP4_23_INFUNC_EN 0
`define DP4_23_OUTFUNC_SEL 0
`define DP4_23_PINCTRL_0_IE 0
`define DP4_23_PINCTRL_0_OD 0
`define DP4_23_PULLEN 0
`define DP4_23_PULLSEL 0
`define DP4_23_pad_y 0
`define DP4_24 0
`define DP4_24_GPIO_OUTPUT_ENABLE 0
`define DP4_24_INFUNC_EN 0
`define DP4_24_OUTFUNC_SEL 0
`define DP4_24_PINCTRL_0_IE 0
`define DP4_24_PINCTRL_0_OD 0
`define DP4_24_PULLEN 0
`define DP4_24_PULLSEL 0
`define DP4_24_pad_y 0
`define DP4_25 0
`define DP4_25_GPIO_OUTPUT_ENABLE 0
`define DP4_25_INFUNC_EN 0
`define DP4_25_OUTFUNC_SEL 0
`define DP4_25_PINCTRL_0_IE 0
`define DP4_25_PINCTRL_0_OD 0
`define DP4_25_PULLEN 0
`define DP4_25_PULLSEL 0
`define DP4_25_pad_y 0
`define DP4_26 0
`define DP4_26_GPIO_OUTPUT_ENABLE 0
`define DP4_26_INFUNC_EN 0
`define DP4_26_OUTFUNC_SEL 0
`define DP4_26_PINCTRL_0_IE 0
`define DP4_26_PINCTRL_0_OD 0
`define DP4_26_PULLEN 0
`define DP4_26_PULLSEL 0
`define DP4_26_pad_y 0
`define DP4_27 0
`define DP4_27_GPIO_OUTPUT_ENABLE 0
`define DP4_27_INFUNC_EN 0
`define DP4_27_OUTFUNC_SEL 0
`define DP4_27_PINCTRL_0_IE 0
`define DP4_27_PINCTRL_0_OD 0
`define DP4_27_PULLEN 0
`define DP4_27_PULLSEL 0
`define DP4_27_pad_y 0
`define DP4_28 0
`define DP4_28_GPIO_OUTPUT_ENABLE 0
`define DP4_28_INFUNC_EN 0
`define DP4_28_OUTFUNC_SEL 0
`define DP4_28_PINCTRL_0_IE 0
`define DP4_28_PINCTRL_0_OD 0
`define DP4_28_PULLEN 0
`define DP4_28_PULLSEL 0
`define DP4_28_pad_y 0
`define DP4_29 0
`define DP4_29_GPIO_OUTPUT_ENABLE 0
`define DP4_29_INFUNC_EN 0
`define DP4_29_OUTFUNC_SEL 0
`define DP4_29_PINCTRL_0_IE 0
`define DP4_29_PINCTRL_0_OD 0
`define DP4_29_PULLEN 0
`define DP4_29_PULLSEL 0
`define DP4_29_pad_y 0
`define DP4_2_GPIO_OUTPUT_ENABLE 0
`define DP4_2_INFUNC_EN 0
`define DP4_2_OUTFUNC_SEL 0
`define DP4_2_PINCTRL_0_IE 0
`define DP4_2_PINCTRL_0_OD 0
`define DP4_2_PULLEN 0
`define DP4_2_PULLSEL 0
`define DP4_2_pad_y 0
`define DP4_3 0
`define DP4_30 0
`define DP4_30_GPIO_OUTPUT_ENABLE 0
`define DP4_30_INFUNC_EN 0
`define DP4_30_OUTFUNC_SEL 0
`define DP4_30_PINCTRL_0_IE 0
`define DP4_30_PINCTRL_0_OD 0
`define DP4_30_PULLEN 0
`define DP4_30_PULLSEL 0
`define DP4_30_pad_y 0
`define DP4_31 0
`define DP4_31_GPIO_OUTPUT_ENABLE 0
`define DP4_31_INFUNC_EN 0
`define DP4_31_OUTFUNC_SEL 0
`define DP4_31_PINCTRL_0_IE 0
`define DP4_31_PINCTRL_0_OD 0
`define DP4_31_PULLEN 0
`define DP4_31_PULLSEL 0
`define DP4_31_pad_y 0
`define DP4_3_GPIO_OUTPUT_ENABLE 0
`define DP4_3_INFUNC_EN 0
`define DP4_3_OUTFUNC_SEL 0
`define DP4_3_PINCTRL_0_IE 0
`define DP4_3_PINCTRL_0_OD 0
`define DP4_3_PULLEN 0
`define DP4_3_PULLSEL 0
`define DP4_3_pad_y 0
`define DP4_4 0
`define DP4_4_GPIO_OUTPUT_ENABLE 0
`define DP4_4_INFUNC_EN 0
`define DP4_4_OUTFUNC_SEL 0
`define DP4_4_PINCTRL_0_IE 0
`define DP4_4_PINCTRL_0_OD 0
`define DP4_4_PULLEN 0
`define DP4_4_PULLSEL 0
`define DP4_4_pad_y 0
`define DP4_5 0
`define DP4_5_GPIO_OUTPUT_ENABLE 0
`define DP4_5_INFUNC_EN 0
`define DP4_5_OUTFUNC_SEL 0
`define DP4_5_PINCTRL_0_IE 0
`define DP4_5_PINCTRL_0_OD 0
`define DP4_5_PULLEN 0
`define DP4_5_PULLSEL 0
`define DP4_5_pad_y 0
`define DP4_6 0
`define DP4_6_GPIO_OUTPUT_ENABLE 0
`define DP4_6_INFUNC_EN 0
`define DP4_6_OUTFUNC_SEL 0
`define DP4_6_PINCTRL_0_IE 0
`define DP4_6_PINCTRL_0_OD 0
`define DP4_6_PULLEN 0
`define DP4_6_PULLSEL 0
`define DP4_6_pad_y 0
`define DP4_7 0
`define DP4_7_GPIO_OUTPUT_ENABLE 0
`define DP4_7_INFUNC_EN 0
`define DP4_7_OUTFUNC_SEL 0
`define DP4_7_PINCTRL_0_IE 0
`define DP4_7_PINCTRL_0_OD 0
`define DP4_7_PULLEN 0
`define DP4_7_PULLSEL 0
`define DP4_7_pad_y 0
`define DP4_8 0
`define DP4_8_GPIO_OUTPUT_ENABLE 0
`define DP4_8_INFUNC_EN 0
`define DP4_8_OUTFUNC_SEL 0
`define DP4_8_PINCTRL_0_IE 0
`define DP4_8_PINCTRL_0_OD 0
`define DP4_8_PULLEN 0
`define DP4_8_PULLSEL 0
`define DP4_8_pad_y 0
`define DP4_9 0
`define DP4_9_GPIO_OUTPUT_ENABLE 0
`define DP4_9_INFUNC_EN 0
`define DP4_9_OUTFUNC_SEL 0
`define DP4_9_PINCTRL_0_IE 0
`define DP4_9_PINCTRL_0_OD 0
`define DP4_9_PULLEN 0
`define DP4_9_PULLSEL 0
`define DP4_9_pad_y 0
`define DP5_0 0
`define DP5_0_GPIO_OUTPUT_ENABLE 0
`define DP5_0_INFUNC_EN 0
`define DP5_0_OUTFUNC_SEL 0
`define DP5_0_PINCTRL_0_IE 0
`define DP5_0_PINCTRL_0_OD 0
`define DP5_0_PULLEN 0
`define DP5_0_PULLSEL 0
`define DP5_0_pad_y 0
`define DP5_1 0
`define DP5_10 0
`define DP5_10_GPIO_OUTPUT_ENABLE 0
`define DP5_10_INFUNC_EN 0
`define DP5_10_OUTFUNC_SEL 0
`define DP5_10_PINCTRL_0_IE 0
`define DP5_10_PINCTRL_0_OD 0
`define DP5_10_PULLEN 0
`define DP5_10_PULLSEL 0
`define DP5_10_pad_y 0
`define DP5_11 0
`define DP5_11_GPIO_OUTPUT_ENABLE 0
`define DP5_11_INFUNC_EN 0
`define DP5_11_OUTFUNC_SEL 0
`define DP5_11_PINCTRL_0_IE 0
`define DP5_11_PINCTRL_0_OD 0
`define DP5_11_PULLEN 0
`define DP5_11_PULLSEL 0
`define DP5_11_pad_y 0
`define DP5_12 0
`define DP5_12_GPIO_OUTPUT_ENABLE 0
`define DP5_12_INFUNC_EN 0
`define DP5_12_OUTFUNC_SEL 0
`define DP5_12_PINCTRL_0_IE 0
`define DP5_12_PINCTRL_0_OD 0
`define DP5_12_PULLEN 0
`define DP5_12_PULLSEL 0
`define DP5_12_pad_y 0
`define DP5_13 0
`define DP5_13_GPIO_OUTPUT_ENABLE 0
`define DP5_13_INFUNC_EN 0
`define DP5_13_OUTFUNC_SEL 0
`define DP5_13_PINCTRL_0_IE 0
`define DP5_13_PINCTRL_0_OD 0
`define DP5_13_PULLEN 0
`define DP5_13_PULLSEL 0
`define DP5_13_pad_y 0
`define DP5_14 0
`define DP5_14_GPIO_OUTPUT_ENABLE 0
`define DP5_14_INFUNC_EN 0
`define DP5_14_OUTFUNC_SEL 0
`define DP5_14_PINCTRL_0_IE 0
`define DP5_14_PINCTRL_0_OD 0
`define DP5_14_PULLEN 0
`define DP5_14_PULLSEL 0
`define DP5_14_pad_y 0
`define DP5_15 0
`define DP5_15_GPIO_OUTPUT_ENABLE 0
`define DP5_15_INFUNC_EN 0
`define DP5_15_OUTFUNC_SEL 0
`define DP5_15_PINCTRL_0_IE 0
`define DP5_15_PINCTRL_0_OD 0
`define DP5_15_PULLEN 0
`define DP5_15_PULLSEL 0
`define DP5_15_pad_y 0
`define DP5_16 0
`define DP5_16_GPIO_OUTPUT_ENABLE 0
`define DP5_16_INFUNC_EN 0
`define DP5_16_OUTFUNC_SEL 0
`define DP5_16_PINCTRL_0_IE 0
`define DP5_16_PINCTRL_0_OD 0
`define DP5_16_PULLEN 0
`define DP5_16_PULLSEL 0
`define DP5_16_pad_y 0
`define DP5_17 0
`define DP5_17_GPIO_OUTPUT_ENABLE 0
`define DP5_17_INFUNC_EN 0
`define DP5_17_OUTFUNC_SEL 0
`define DP5_17_PINCTRL_0_IE 0
`define DP5_17_PINCTRL_0_OD 0
`define DP5_17_PULLEN 0
`define DP5_17_PULLSEL 0
`define DP5_17_pad_y 0
`define DP5_18 0
`define DP5_18_GPIO_OUTPUT_ENABLE 0
`define DP5_18_INFUNC_EN 0
`define DP5_18_OUTFUNC_SEL 0
`define DP5_18_PINCTRL_0_IE 0
`define DP5_18_PINCTRL_0_OD 0
`define DP5_18_PULLEN 0
`define DP5_18_PULLSEL 0
`define DP5_18_pad_y 0
`define DP5_19 0
`define DP5_19_GPIO_OUTPUT_ENABLE 0
`define DP5_19_INFUNC_EN 0
`define DP5_19_OUTFUNC_SEL 0
`define DP5_19_PINCTRL_0_IE 0
`define DP5_19_PINCTRL_0_OD 0
`define DP5_19_PULLEN 0
`define DP5_19_PULLSEL 0
`define DP5_19_pad_y 0
`define DP5_1_GPIO_OUTPUT_ENABLE 0
`define DP5_1_INFUNC_EN 0
`define DP5_1_OUTFUNC_SEL 0
`define DP5_1_PINCTRL_0_IE 0
`define DP5_1_PINCTRL_0_OD 0
`define DP5_1_PULLEN 0
`define DP5_1_PULLSEL 0
`define DP5_1_pad_y 0
`define DP5_2 0
`define DP5_20 0
`define DP5_20_GPIO_OUTPUT_ENABLE 0
`define DP5_20_INFUNC_EN 0
`define DP5_20_OUTFUNC_SEL 0
`define DP5_20_PINCTRL_0_IE 0
`define DP5_20_PINCTRL_0_OD 0
`define DP5_20_PULLEN 0
`define DP5_20_PULLSEL 0
`define DP5_20_pad_y 0
`define DP5_21 0
`define DP5_21_GPIO_OUTPUT_ENABLE 0
`define DP5_21_INFUNC_EN 0
`define DP5_21_OUTFUNC_SEL 0
`define DP5_21_PINCTRL_0_IE 0
`define DP5_21_PINCTRL_0_OD 0
`define DP5_21_PULLEN 0
`define DP5_21_PULLSEL 0
`define DP5_21_pad_y 0
`define DP5_22 0
`define DP5_22_GPIO_OUTPUT_ENABLE 0
`define DP5_22_INFUNC_EN 0
`define DP5_22_OUTFUNC_SEL 0
`define DP5_22_PINCTRL_0_IE 0
`define DP5_22_PINCTRL_0_OD 0
`define DP5_22_PULLEN 0
`define DP5_22_PULLSEL 0
`define DP5_22_pad_y 0
`define DP5_23 0
`define DP5_23_GPIO_OUTPUT_ENABLE 0
`define DP5_23_INFUNC_EN 0
`define DP5_23_OUTFUNC_SEL 0
`define DP5_23_PINCTRL_0_IE 0
`define DP5_23_PINCTRL_0_OD 0
`define DP5_23_PULLEN 0
`define DP5_23_PULLSEL 0
`define DP5_23_pad_y 0
`define DP5_24 0
`define DP5_24_GPIO_OUTPUT_ENABLE 0
`define DP5_24_INFUNC_EN 0
`define DP5_24_OUTFUNC_SEL 0
`define DP5_24_PINCTRL_0_IE 0
`define DP5_24_PINCTRL_0_OD 0
`define DP5_24_PULLEN 0
`define DP5_24_PULLSEL 0
`define DP5_24_pad_y 0
`define DP5_25 0
`define DP5_25_GPIO_OUTPUT_ENABLE 0
`define DP5_25_INFUNC_EN 0
`define DP5_25_OUTFUNC_SEL 0
`define DP5_25_PINCTRL_0_IE 0
`define DP5_25_PINCTRL_0_OD 0
`define DP5_25_PULLEN 0
`define DP5_25_PULLSEL 0
`define DP5_25_pad_y 0
`define DP5_26 0
`define DP5_26_GPIO_OUTPUT_ENABLE 0
`define DP5_26_INFUNC_EN 0
`define DP5_26_OUTFUNC_SEL 0
`define DP5_26_PINCTRL_0_IE 0
`define DP5_26_PINCTRL_0_OD 0
`define DP5_26_PULLEN 0
`define DP5_26_PULLSEL 0
`define DP5_26_pad_y 0
`define DP5_27 0
`define DP5_27_GPIO_OUTPUT_ENABLE 0
`define DP5_27_INFUNC_EN 0
`define DP5_27_OUTFUNC_SEL 0
`define DP5_27_PINCTRL_0_IE 0
`define DP5_27_PINCTRL_0_OD 0
`define DP5_27_PULLEN 0
`define DP5_27_PULLSEL 0
`define DP5_27_pad_y 0
`define DP5_28 0
`define DP5_28_GPIO_OUTPUT_ENABLE 0
`define DP5_28_INFUNC_EN 0
`define DP5_28_OUTFUNC_SEL 0
`define DP5_28_PINCTRL_0_IE 0
`define DP5_28_PINCTRL_0_OD 0
`define DP5_28_PULLEN 0
`define DP5_28_PULLSEL 0
`define DP5_28_pad_y 0
`define DP5_29 0
`define DP5_29_GPIO_OUTPUT_ENABLE 0
`define DP5_29_INFUNC_EN 0
`define DP5_29_OUTFUNC_SEL 0
`define DP5_29_PINCTRL_0_IE 0
`define DP5_29_PINCTRL_0_OD 0
`define DP5_29_PULLEN 0
`define DP5_29_PULLSEL 0
`define DP5_29_pad_y 0
`define DP5_2_GPIO_OUTPUT_ENABLE 0
`define DP5_2_INFUNC_EN 0
`define DP5_2_OUTFUNC_SEL 0
`define DP5_2_PINCTRL_0_IE 0
`define DP5_2_PINCTRL_0_OD 0
`define DP5_2_PULLEN 0
`define DP5_2_PULLSEL 0
`define DP5_2_pad_y 0
`define DP5_3 0
`define DP5_30 0
`define DP5_30_GPIO_OUTPUT_ENABLE 0
`define DP5_30_INFUNC_EN 0
`define DP5_30_OUTFUNC_SEL 0
`define DP5_30_PINCTRL_0_IE 0
`define DP5_30_PINCTRL_0_OD 0
`define DP5_30_PULLEN 0
`define DP5_30_PULLSEL 0
`define DP5_30_pad_y 0
`define DP5_31 0
`define DP5_31_GPIO_OUTPUT_ENABLE 0
`define DP5_31_INFUNC_EN 0
`define DP5_31_OUTFUNC_SEL 0
`define DP5_31_PINCTRL_0_IE 0
`define DP5_31_PINCTRL_0_OD 0
`define DP5_31_PULLEN 0
`define DP5_31_PULLSEL 0
`define DP5_31_pad_y 0
`define DP5_3_GPIO_OUTPUT_ENABLE 0
`define DP5_3_INFUNC_EN 0
`define DP5_3_OUTFUNC_SEL 0
`define DP5_3_PINCTRL_0_IE 0
`define DP5_3_PINCTRL_0_OD 0
`define DP5_3_PULLEN 0
`define DP5_3_PULLSEL 0
`define DP5_3_pad_y 0
`define DP5_4 0
`define DP5_4_GPIO_OUTPUT_ENABLE 0
`define DP5_4_INFUNC_EN 0
`define DP5_4_OUTFUNC_SEL 0
`define DP5_4_PINCTRL_0_IE 0
`define DP5_4_PINCTRL_0_OD 0
`define DP5_4_PULLEN 0
`define DP5_4_PULLSEL 0
`define DP5_4_pad_y 0
`define DP5_5 0
`define DP5_5_GPIO_OUTPUT_ENABLE 0
`define DP5_5_INFUNC_EN 0
`define DP5_5_OUTFUNC_SEL 0
`define DP5_5_PINCTRL_0_IE 0
`define DP5_5_PINCTRL_0_OD 0
`define DP5_5_PULLEN 0
`define DP5_5_PULLSEL 0
`define DP5_5_pad_y 0
`define DP5_6 0
`define DP5_6_GPIO_OUTPUT_ENABLE 0
`define DP5_6_INFUNC_EN 0
`define DP5_6_OUTFUNC_SEL 0
`define DP5_6_PINCTRL_0_IE 0
`define DP5_6_PINCTRL_0_OD 0
`define DP5_6_PULLEN 0
`define DP5_6_PULLSEL 0
`define DP5_6_pad_y 0
`define DP5_7 0
`define DP5_7_GPIO_OUTPUT_ENABLE 0
`define DP5_7_INFUNC_EN 0
`define DP5_7_OUTFUNC_SEL 0
`define DP5_7_PINCTRL_0_IE 0
`define DP5_7_PINCTRL_0_OD 0
`define DP5_7_PULLEN 0
`define DP5_7_PULLSEL 0
`define DP5_7_pad_y 0
`define DP5_8 0
`define DP5_8_GPIO_OUTPUT_ENABLE 0
`define DP5_8_INFUNC_EN 0
`define DP5_8_OUTFUNC_SEL 0
`define DP5_8_PINCTRL_0_IE 0
`define DP5_8_PINCTRL_0_OD 0
`define DP5_8_PULLEN 0
`define DP5_8_PULLSEL 0
`define DP5_8_pad_y 0
`define DP5_9 0
`define DP5_9_GPIO_OUTPUT_ENABLE 0
`define DP5_9_INFUNC_EN 0
`define DP5_9_OUTFUNC_SEL 0
`define DP5_9_PINCTRL_0_IE 0
`define DP5_9_PINCTRL_0_OD 0
`define DP5_9_PULLEN 0
`define DP5_9_PULLSEL 0
`define DP5_9_pad_y 0
`define DP6_0 0
`define DP6_0_GPIO_OUTPUT_ENABLE 0
`define DP6_0_INFUNC_EN 0
`define DP6_0_OUTFUNC_SEL 0
`define DP6_0_PINCTRL_0_IE 0
`define DP6_0_PINCTRL_0_OD 0
`define DP6_0_PULLEN 0
`define DP6_0_PULLSEL 0
`define DP6_0_pad_y 0
`define DP6_1 0
`define DP6_10 0
`define DP6_10_GPIO_OUTPUT_ENABLE 0
`define DP6_10_INFUNC_EN 0
`define DP6_10_OUTFUNC_SEL 0
`define DP6_10_PINCTRL_0_IE 0
`define DP6_10_PINCTRL_0_OD 0
`define DP6_10_PULLEN 0
`define DP6_10_PULLSEL 0
`define DP6_10_pad_y 0
`define DP6_11 0
`define DP6_11_GPIO_OUTPUT_ENABLE 0
`define DP6_11_INFUNC_EN 0
`define DP6_11_OUTFUNC_SEL 0
`define DP6_11_PINCTRL_0_IE 0
`define DP6_11_PINCTRL_0_OD 0
`define DP6_11_PULLEN 0
`define DP6_11_PULLSEL 0
`define DP6_11_pad_y 0
`define DP6_12 0
`define DP6_12_GPIO_OUTPUT_ENABLE 0
`define DP6_12_INFUNC_EN 0
`define DP6_12_OUTFUNC_SEL 0
`define DP6_12_PINCTRL_0_IE 0
`define DP6_12_PINCTRL_0_OD 0
`define DP6_12_PULLEN 0
`define DP6_12_PULLSEL 0
`define DP6_12_pad_y 0
`define DP6_13 0
`define DP6_13_GPIO_OUTPUT_ENABLE 0
`define DP6_13_INFUNC_EN 0
`define DP6_13_OUTFUNC_SEL 0
`define DP6_13_PINCTRL_0_IE 0
`define DP6_13_PINCTRL_0_OD 0
`define DP6_13_PULLEN 0
`define DP6_13_PULLSEL 0
`define DP6_13_pad_y 0
`define DP6_14 0
`define DP6_14_GPIO_OUTPUT_ENABLE 0
`define DP6_14_INFUNC_EN 0
`define DP6_14_OUTFUNC_SEL 0
`define DP6_14_PINCTRL_0_IE 0
`define DP6_14_PINCTRL_0_OD 0
`define DP6_14_PULLEN 0
`define DP6_14_PULLSEL 0
`define DP6_14_pad_y 0
`define DP6_15 0
`define DP6_15_GPIO_OUTPUT_ENABLE 0
`define DP6_15_INFUNC_EN 0
`define DP6_15_OUTFUNC_SEL 0
`define DP6_15_PINCTRL_0_IE 0
`define DP6_15_PINCTRL_0_OD 0
`define DP6_15_PULLEN 0
`define DP6_15_PULLSEL 0
`define DP6_15_pad_y 0
`define DP6_16 0
`define DP6_16_GPIO_OUTPUT_ENABLE 0
`define DP6_16_INFUNC_EN 0
`define DP6_16_OUTFUNC_SEL 0
`define DP6_16_PINCTRL_0_IE 0
`define DP6_16_PINCTRL_0_OD 0
`define DP6_16_PULLEN 0
`define DP6_16_PULLSEL 0
`define DP6_16_pad_y 0
`define DP6_17 0
`define DP6_17_GPIO_OUTPUT_ENABLE 0
`define DP6_17_INFUNC_EN 0
`define DP6_17_OUTFUNC_SEL 0
`define DP6_17_PINCTRL_0_IE 0
`define DP6_17_PINCTRL_0_OD 0
`define DP6_17_PULLEN 0
`define DP6_17_PULLSEL 0
`define DP6_17_pad_y 0
`define DP6_18 0
`define DP6_18_GPIO_OUTPUT_ENABLE 0
`define DP6_18_INFUNC_EN 0
`define DP6_18_OUTFUNC_SEL 0
`define DP6_18_PINCTRL_0_IE 0
`define DP6_18_PINCTRL_0_OD 0
`define DP6_18_PULLEN 0
`define DP6_18_PULLSEL 0
`define DP6_18_pad_y 0
`define DP6_19 0
`define DP6_19_GPIO_OUTPUT_ENABLE 0
`define DP6_19_INFUNC_EN 0
`define DP6_19_OUTFUNC_SEL 0
`define DP6_19_PINCTRL_0_IE 0
`define DP6_19_PINCTRL_0_OD 0
`define DP6_19_PULLEN 0
`define DP6_19_PULLSEL 0
`define DP6_19_pad_y 0
`define DP6_1_GPIO_OUTPUT_ENABLE 0
`define DP6_1_INFUNC_EN 0
`define DP6_1_OUTFUNC_SEL 0
`define DP6_1_PINCTRL_0_IE 0
`define DP6_1_PINCTRL_0_OD 0
`define DP6_1_PULLEN 0
`define DP6_1_PULLSEL 0
`define DP6_1_pad_y 0
`define DP6_2 0
`define DP6_20 0
`define DP6_20_GPIO_OUTPUT_ENABLE 0
`define DP6_20_INFUNC_EN 0
`define DP6_20_OUTFUNC_SEL 0
`define DP6_20_PINCTRL_0_IE 0
`define DP6_20_PINCTRL_0_OD 0
`define DP6_20_PULLEN 0
`define DP6_20_PULLSEL 0
`define DP6_20_pad_y 0
`define DP6_21 0
`define DP6_21_GPIO_OUTPUT_ENABLE 0
`define DP6_21_INFUNC_EN 0
`define DP6_21_OUTFUNC_SEL 0
`define DP6_21_PINCTRL_0_IE 0
`define DP6_21_PINCTRL_0_OD 0
`define DP6_21_PULLEN 0
`define DP6_21_PULLSEL 0
`define DP6_21_pad_y 0
`define DP6_22 0
`define DP6_22_GPIO_OUTPUT_ENABLE 0
`define DP6_22_INFUNC_EN 0
`define DP6_22_OUTFUNC_SEL 0
`define DP6_22_PINCTRL_0_IE 0
`define DP6_22_PINCTRL_0_OD 0
`define DP6_22_PULLEN 0
`define DP6_22_PULLSEL 0
`define DP6_22_pad_y 0
`define DP6_23 0
`define DP6_23_GPIO_OUTPUT_ENABLE 0
`define DP6_23_INFUNC_EN 0
`define DP6_23_OUTFUNC_SEL 0
`define DP6_23_PINCTRL_0_IE 0
`define DP6_23_PINCTRL_0_OD 0
`define DP6_23_PULLEN 0
`define DP6_23_PULLSEL 0
`define DP6_23_pad_y 0
`define DP6_24 0
`define DP6_24_GPIO_OUTPUT_ENABLE 0
`define DP6_24_INFUNC_EN 0
`define DP6_24_OUTFUNC_SEL 0
`define DP6_24_PINCTRL_0_IE 0
`define DP6_24_PINCTRL_0_OD 0
`define DP6_24_PULLEN 0
`define DP6_24_PULLSEL 0
`define DP6_24_pad_y 0
`define DP6_25 0
`define DP6_25_GPIO_OUTPUT_ENABLE 0
`define DP6_25_INFUNC_EN 0
`define DP6_25_OUTFUNC_SEL 0
`define DP6_25_PINCTRL_0_IE 0
`define DP6_25_PINCTRL_0_OD 0
`define DP6_25_PULLEN 0
`define DP6_25_PULLSEL 0
`define DP6_25_pad_y 0
`define DP6_26 0
`define DP6_26_GPIO_OUTPUT_ENABLE 0
`define DP6_26_INFUNC_EN 0
`define DP6_26_OUTFUNC_SEL 0
`define DP6_26_PINCTRL_0_IE 0
`define DP6_26_PINCTRL_0_OD 0
`define DP6_26_PULLEN 0
`define DP6_26_PULLSEL 0
`define DP6_26_pad_y 0
`define DP6_27 0
`define DP6_27_GPIO_OUTPUT_ENABLE 0
`define DP6_27_INFUNC_EN 0
`define DP6_27_OUTFUNC_SEL 0
`define DP6_27_PINCTRL_0_IE 0
`define DP6_27_PINCTRL_0_OD 0
`define DP6_27_PULLEN 0
`define DP6_27_PULLSEL 0
`define DP6_27_pad_y 0
`define DP6_2_GPIO_OUTPUT_ENABLE 0
`define DP6_2_INFUNC_EN 0
`define DP6_2_OUTFUNC_SEL 0
`define DP6_2_PINCTRL_0_IE 0
`define DP6_2_PINCTRL_0_OD 0
`define DP6_2_PULLEN 0
`define DP6_2_PULLSEL 0
`define DP6_2_pad_y 0
`define DP6_3 0
`define DP6_3_GPIO_OUTPUT_ENABLE 0
`define DP6_3_INFUNC_EN 0
`define DP6_3_OUTFUNC_SEL 0
`define DP6_3_PINCTRL_0_IE 0
`define DP6_3_PINCTRL_0_OD 0
`define DP6_3_PULLEN 0
`define DP6_3_PULLSEL 0
`define DP6_3_pad_y 0
`define DP6_4 0
`define DP6_4_GPIO_OUTPUT_ENABLE 0
`define DP6_4_INFUNC_EN 0
`define DP6_4_OUTFUNC_SEL 0
`define DP6_4_PINCTRL_0_IE 0
`define DP6_4_PINCTRL_0_OD 0
`define DP6_4_PULLEN 0
`define DP6_4_PULLSEL 0
`define DP6_4_pad_y 0
`define DP6_5 0
`define DP6_5_GPIO_OUTPUT_ENABLE 0
`define DP6_5_INFUNC_EN 0
`define DP6_5_OUTFUNC_SEL 0
`define DP6_5_PINCTRL_0_IE 0
`define DP6_5_PINCTRL_0_OD 0
`define DP6_5_PULLEN 0
`define DP6_5_PULLSEL 0
`define DP6_5_pad_y 0
`define DP6_6 0
`define DP6_6_GPIO_OUTPUT_ENABLE 0
`define DP6_6_INFUNC_EN 0
`define DP6_6_OUTFUNC_SEL 0
`define DP6_6_PINCTRL_0_IE 0
`define DP6_6_PINCTRL_0_OD 0
`define DP6_6_PULLEN 0
`define DP6_6_PULLSEL 0
`define DP6_6_pad_y 0
`define DP6_7 0
`define DP6_7_GPIO_OUTPUT_ENABLE 0
`define DP6_7_INFUNC_EN 0
`define DP6_7_OUTFUNC_SEL 0
`define DP6_7_PINCTRL_0_IE 0
`define DP6_7_PINCTRL_0_OD 0
`define DP6_7_PULLEN 0
`define DP6_7_PULLSEL 0
`define DP6_7_pad_y 0
`define DP6_8 0
`define DP6_8_GPIO_OUTPUT_ENABLE 0
`define DP6_8_INFUNC_EN 0
`define DP6_8_OUTFUNC_SEL 0
`define DP6_8_PINCTRL_0_IE 0
`define DP6_8_PINCTRL_0_OD 0
`define DP6_8_PULLEN 0
`define DP6_8_PULLSEL 0
`define DP6_8_pad_y 0
`define DP6_9 0
`define DP6_9_GPIO_OUTPUT_ENABLE 0
`define DP6_9_INFUNC_EN 0
`define DP6_9_OUTFUNC_SEL 0
`define DP6_9_PINCTRL_0_IE 0
`define DP6_9_PINCTRL_0_OD 0
`define DP6_9_PULLEN 0
`define DP6_9_PULLSEL 0
`define DP6_9_pad_y 0
`define DP7_0 0
`define DP7_0_GPIO_OUTPUT_ENABLE 0
`define DP7_0_INFUNC_EN 0
`define DP7_0_OUTFUNC_SEL 0
`define DP7_0_PINCTRL_0_IE 0
`define DP7_0_PINCTRL_0_OD 0
`define DP7_0_PULLEN 0
`define DP7_0_PULLSEL 0
`define DP7_0_pad_y 0
`define DP7_1 0
`define DP7_10 0
`define DP7_10_GPIO_OUTPUT_ENABLE 0
`define DP7_10_INFUNC_EN 0
`define DP7_10_OUTFUNC_SEL 0
`define DP7_10_PINCTRL_0_IE 0
`define DP7_10_PINCTRL_0_OD 0
`define DP7_10_PULLEN 0
`define DP7_10_PULLSEL 0
`define DP7_10_pad_y 0
`define DP7_11 0
`define DP7_11_GPIO_OUTPUT_ENABLE 0
`define DP7_11_INFUNC_EN 0
`define DP7_11_OUTFUNC_SEL 0
`define DP7_11_PINCTRL_0_IE 0
`define DP7_11_PINCTRL_0_OD 0
`define DP7_11_PULLEN 0
`define DP7_11_PULLSEL 0
`define DP7_11_pad_y 0
`define DP7_12 0
`define DP7_12_GPIO_OUTPUT_ENABLE 0
`define DP7_12_INFUNC_EN 0
`define DP7_12_OUTFUNC_SEL 0
`define DP7_12_PINCTRL_0_IE 0
`define DP7_12_PINCTRL_0_OD 0
`define DP7_12_PULLEN 0
`define DP7_12_PULLSEL 0
`define DP7_12_pad_y 0
`define DP7_13 0
`define DP7_13_GPIO_OUTPUT_ENABLE 0
`define DP7_13_INFUNC_EN 0
`define DP7_13_OUTFUNC_SEL 0
`define DP7_13_PINCTRL_0_IE 0
`define DP7_13_PINCTRL_0_OD 0
`define DP7_13_PULLEN 0
`define DP7_13_PULLSEL 0
`define DP7_13_pad_y 0
`define DP7_14 0
`define DP7_14_GPIO_OUTPUT_ENABLE 0
`define DP7_14_INFUNC_EN 0
`define DP7_14_OUTFUNC_SEL 0
`define DP7_14_PINCTRL_0_IE 0
`define DP7_14_PINCTRL_0_OD 0
`define DP7_14_PULLEN 0
`define DP7_14_PULLSEL 0
`define DP7_14_pad_y 0
`define DP7_15 0
`define DP7_15_GPIO_OUTPUT_ENABLE 0
`define DP7_15_INFUNC_EN 0
`define DP7_15_OUTFUNC_SEL 0
`define DP7_15_PINCTRL_0_IE 0
`define DP7_15_PINCTRL_0_OD 0
`define DP7_15_PULLEN 0
`define DP7_15_PULLSEL 0
`define DP7_15_pad_y 0
`define DP7_1_GPIO_OUTPUT_ENABLE 0
`define DP7_1_INFUNC_EN 0
`define DP7_1_OUTFUNC_SEL 0
`define DP7_1_PINCTRL_0_IE 0
`define DP7_1_PINCTRL_0_OD 0
`define DP7_1_PULLEN 0
`define DP7_1_PULLSEL 0
`define DP7_1_pad_y 0
`define DP7_2 0
`define DP7_2_GPIO_OUTPUT_ENABLE 0
`define DP7_2_INFUNC_EN 0
`define DP7_2_OUTFUNC_SEL 0
`define DP7_2_PINCTRL_0_IE 0
`define DP7_2_PINCTRL_0_OD 0
`define DP7_2_PULLEN 0
`define DP7_2_PULLSEL 0
`define DP7_2_pad_y 0
`define DP7_3 0
`define DP7_3_GPIO_OUTPUT_ENABLE 0
`define DP7_3_INFUNC_EN 0
`define DP7_3_OUTFUNC_SEL 0
`define DP7_3_PINCTRL_0_IE 0
`define DP7_3_PINCTRL_0_OD 0
`define DP7_3_PULLEN 0
`define DP7_3_PULLSEL 0
`define DP7_3_pad_y 0
`define DP7_4 0
`define DP7_4_GPIO_OUTPUT_ENABLE 0
`define DP7_4_INFUNC_EN 0
`define DP7_4_OUTFUNC_SEL 0
`define DP7_4_PINCTRL_0_IE 0
`define DP7_4_PINCTRL_0_OD 0
`define DP7_4_PULLEN 0
`define DP7_4_PULLSEL 0
`define DP7_4_pad_y 0
`define DP7_5 0
`define DP7_5_GPIO_OUTPUT_ENABLE 0
`define DP7_5_INFUNC_EN 0
`define DP7_5_OUTFUNC_SEL 0
`define DP7_5_PINCTRL_0_IE 0
`define DP7_5_PINCTRL_0_OD 0
`define DP7_5_PULLEN 0
`define DP7_5_PULLSEL 0
`define DP7_5_pad_y 0
`define DP7_6 0
`define DP7_6_GPIO_OUTPUT_ENABLE 0
`define DP7_6_INFUNC_EN 0
`define DP7_6_OUTFUNC_SEL 0
`define DP7_6_PINCTRL_0_IE 0
`define DP7_6_PINCTRL_0_OD 0
`define DP7_6_PULLEN 0
`define DP7_6_PULLSEL 0
`define DP7_6_pad_y 0
`define DP7_7 0
`define DP7_7_GPIO_OUTPUT_ENABLE 0
`define DP7_7_INFUNC_EN 0
`define DP7_7_OUTFUNC_SEL 0
`define DP7_7_PINCTRL_0_IE 0
`define DP7_7_PINCTRL_0_OD 0
`define DP7_7_PULLEN 0
`define DP7_7_PULLSEL 0
`define DP7_7_pad_y 0
`define DP7_8 0
`define DP7_8_GPIO_OUTPUT_ENABLE 0
`define DP7_8_INFUNC_EN 0
`define DP7_8_OUTFUNC_SEL 0
`define DP7_8_PINCTRL_0_IE 0
`define DP7_8_PINCTRL_0_OD 0
`define DP7_8_PULLEN 0
`define DP7_8_PULLSEL 0
`define DP7_8_pad_y 0
`define DP7_9 0
`define DP7_9_GPIO_OUTPUT_ENABLE 0
`define DP7_9_INFUNC_EN 0
`define DP7_9_OUTFUNC_SEL 0
`define DP7_9_PINCTRL_0_IE 0
`define DP7_9_PINCTRL_0_OD 0
`define DP7_9_PULLEN 0
`define DP7_9_PULLSEL 0
`define DP7_9_pad_y 0
`define EPWM0A_IN 0
`define EPWM0A_OE 0
`define EPWM0A_OUT 0
`define EPWM0B_IN 0
`define EPWM0B_OE 0
`define EPWM0B_OUT 0
`define EPWM10A_IN 0
`define EPWM10A_OE 0
`define EPWM10A_OUT 0
`define EPWM10B_IN 0
`define EPWM10B_OE 0
`define EPWM10B_OUT 0
`define EPWM11A_IN 0
`define EPWM11A_OE 0
`define EPWM11A_OUT 0
`define EPWM11B_IN 0
`define EPWM11B_OE 0
`define EPWM11B_OUT 0
`define EPWM12A_IN 0
`define EPWM12A_OE 0
`define EPWM12A_OUT 0
`define EPWM12B_IN 0
`define EPWM12B_OE 0
`define EPWM12B_OUT 0
`define EPWM13A_IN 0
`define EPWM13A_OE 0
`define EPWM13A_OUT 0
`define EPWM13B_IN 0
`define EPWM13B_OE 0
`define EPWM13B_OUT 0
`define EPWM14A_IN 0
`define EPWM14A_OE 0
`define EPWM14A_OUT 0
`define EPWM14B_IN 0
`define EPWM14B_OE 0
`define EPWM14B_OUT 0
`define EPWM15A_IN 0
`define EPWM15A_OE 0
`define EPWM15A_OUT 0
`define EPWM15B_IN 0
`define EPWM15B_OE 0
`define EPWM15B_OUT 0
`define EPWM16A_IN 0
`define EPWM16A_OE 0
`define EPWM16A_OUT 0
`define EPWM16B_IN 0
`define EPWM16B_OE 0
`define EPWM16B_OUT 0
`define EPWM17A_IN 0
`define EPWM17A_OE 0
`define EPWM17A_OUT 0
`define EPWM17B_IN 0
`define EPWM17B_OE 0
`define EPWM17B_OUT 0
`define EPWM18A_IN 0
`define EPWM18A_OE 0
`define EPWM18A_OUT 0
`define EPWM18B_IN 0
`define EPWM18B_OE 0
`define EPWM18B_OUT 0
`define EPWM19A_IN 0
`define EPWM19A_OE 0
`define EPWM19A_OUT 0
`define EPWM19B_IN 0
`define EPWM19B_OE 0
`define EPWM19B_OUT 0
`define EPWM1A_IN 0
`define EPWM1A_OE 0
`define EPWM1A_OUT 0
`define EPWM1B_IN 0
`define EPWM1B_OE 0
`define EPWM1B_OUT 0
`define EPWM20A_IN 0
`define EPWM20A_OE 0
`define EPWM20A_OUT 0
`define EPWM20B_IN 0
`define EPWM20B_OE 0
`define EPWM20B_OUT 0
`define EPWM21A_IN 0
`define EPWM21A_OE 0
`define EPWM21A_OUT 0
`define EPWM21B_IN 0
`define EPWM21B_OE 0
`define EPWM21B_OUT 0
`define EPWM22A_IN 0
`define EPWM22A_OE 0
`define EPWM22A_OUT 0
`define EPWM22B_IN 0
`define EPWM22B_OE 0
`define EPWM22B_OUT 0
`define EPWM23A_IN 0
`define EPWM23A_OE 0
`define EPWM23A_OUT 0
`define EPWM23B_IN 0
`define EPWM23B_OE 0
`define EPWM23B_OUT 0
`define EPWM24A_IN 0
`define EPWM24A_OE 0
`define EPWM24A_OUT 0
`define EPWM24B_IN 0
`define EPWM24B_OE 0
`define EPWM24B_OUT 0
`define EPWM25A_IN 0
`define EPWM25A_OE 0
`define EPWM25A_OUT 0
`define EPWM25B_IN 0
`define EPWM25B_OE 0
`define EPWM25B_OUT 0
`define EPWM26A_IN 0
`define EPWM26A_OE 0
`define EPWM26A_OUT 0
`define EPWM26B_IN 0
`define EPWM26B_OE 0
`define EPWM26B_OUT 0
`define EPWM27A_IN 0
`define EPWM27A_OE 0
`define EPWM27A_OUT 0
`define EPWM27B_IN 0
`define EPWM27B_OE 0
`define EPWM27B_OUT 0
`define EPWM28A_IN 0
`define EPWM28A_OE 0
`define EPWM28A_OUT 0
`define EPWM28B_IN 0
`define EPWM28B_OE 0
`define EPWM28B_OUT 0
`define EPWM29A_IN 0
`define EPWM29A_OE 0
`define EPWM29A_OUT 0
`define EPWM29B_IN 0
`define EPWM29B_OE 0
`define EPWM29B_OUT 0
`define EPWM2A_IN 0
`define EPWM2A_OE 0
`define EPWM2A_OUT 0
`define EPWM2B_IN 0
`define EPWM2B_OE 0
`define EPWM2B_OUT 0
`define EPWM30A_IN 0
`define EPWM30A_OE 0
`define EPWM30A_OUT 0
`define EPWM30B_IN 0
`define EPWM30B_OE 0
`define EPWM30B_OUT 0
`define EPWM31A_IN 0
`define EPWM31A_OE 0
`define EPWM31A_OUT 0
`define EPWM31B_IN 0
`define EPWM31B_OE 0
`define EPWM31B_OUT 0
`define EPWM3A_IN 0
`define EPWM3A_OE 0
`define EPWM3A_OUT 0
`define EPWM3B_IN 0
`define EPWM3B_OE 0
`define EPWM3B_OUT 0
`define EPWM4A_IN 0
`define EPWM4A_OE 0
`define EPWM4A_OUT 0
`define EPWM4B_IN 0
`define EPWM4B_OE 0
`define EPWM4B_OUT 0
`define EPWM5A_IN 0
`define EPWM5A_OE 0
`define EPWM5A_OUT 0
`define EPWM5B_IN 0
`define EPWM5B_OE 0
`define EPWM5B_OUT 0
`define EPWM6A_IN 0
`define EPWM6A_OE 0
`define EPWM6A_OUT 0
`define EPWM6B_IN 0
`define EPWM6B_OE 0
`define EPWM6B_OUT 0
`define EPWM7A_IN 0
`define EPWM7A_OE 0
`define EPWM7A_OUT 0
`define EPWM7B_IN 0
`define EPWM7B_OE 0
`define EPWM7B_OUT 0
`define EPWM8A_IN 0
`define EPWM8A_OE 0
`define EPWM8A_OUT 0
`define EPWM8B_IN 0
`define EPWM8B_OE 0
`define EPWM8B_OUT 0
`define EPWM9A_IN 0
`define EPWM9A_OE 0
`define EPWM9A_OUT 0
`define EPWM9B_IN 0
`define EPWM9B_OE 0
`define EPWM9B_OUT 0
`define EPWMSYNCO_IN 0
`define EPWMSYNCO_OE 0
`define EPWMSYNCO_OUT 0
`define EXTCLK_IN 0
`define FSI0RXCLK_IN 0
`define FSI0RXCLK_OE 0
`define FSI0RXCLK_OUT 0
`define FSI0RXD0_IN 0
`define FSI0RXD0_OE 0
`define FSI0RXD0_OUT 0
`define FSI0RXD1_IN 0
`define FSI0RXD1_OE 0
`define FSI0RXD1_OUT 0
`define FSI0TXCLK_IN 0
`define FSI0TXCLK_OE 0
`define FSI0TXCLK_OUT 0
`define FSI0TXD0_IN 0
`define FSI0TXD0_OE 0
`define FSI0TXD0_OUT 0
`define FSI0TXD1_IN 0
`define FSI0TXD1_OE 0
`define FSI0TXD1_OUT 0
`define FSI1RXCLK_IN 0
`define FSI1RXCLK_OE 0
`define FSI1RXCLK_OUT 0
`define FSI1RXD0_IN 0
`define FSI1RXD0_OE 0
`define FSI1RXD0_OUT 0
`define FSI1RXD1_IN 0
`define FSI1RXD1_OE 0
`define FSI1RXD1_OUT 0
`define FSI1TXCLK_IN 0
`define FSI1TXCLK_OE 0
`define FSI1TXCLK_OUT 0
`define FSI1TXD0_IN 0
`define FSI1TXD0_OE 0
`define FSI1TXD0_OUT 0
`define FSI1TXD1_IN 0
`define FSI1TXD1_OE 0
`define FSI1TXD1_OUT 0
`define FSI2RXCLK_IN 0
`define FSI2RXCLK_OE 0
`define FSI2RXCLK_OUT 0
`define FSI2RXD0_IN 0
`define FSI2RXD0_OE 0
`define FSI2RXD0_OUT 0
`define FSI2RXD1_IN 0
`define FSI2RXD1_OE 0
`define FSI2RXD1_OUT 0
`define FSI2TXCLK_IN 0
`define FSI2TXCLK_OE 0
`define FSI2TXCLK_OUT 0
`define FSI2TXD0_IN 0
`define FSI2TXD0_OE 0
`define FSI2TXD0_OUT 0
`define FSI2TXD1_IN 0
`define FSI2TXD1_OE 0
`define FSI2TXD1_OUT 0
`define FSI3RXCLK_IN 0
`define FSI3RXCLK_OE 0
`define FSI3RXCLK_OUT 0
`define FSI3RXD0_IN 0
`define FSI3RXD0_OE 0
`define FSI3RXD0_OUT 0
`define FSI3RXD1_IN 0
`define FSI3RXD1_OE 0
`define FSI3RXD1_OUT 0
`define FSI3TXCLK_IN 0
`define FSI3TXCLK_OE 0
`define FSI3TXCLK_OUT 0
`define FSI3TXD0_IN 0
`define FSI3TXD0_OE 0
`define FSI3TXD0_OUT 0
`define FSI3TXD1_IN 0
`define FSI3TXD1_OE 0
`define FSI3TXD1_OUT 0
`define FSI4RXCLK_IN 0
`define FSI4RXCLK_OE 0
`define FSI4RXCLK_OUT 0
`define FSI4RXD0_IN 0
`define FSI4RXD0_OE 0
`define FSI4RXD0_OUT 0
`define FSI4RXD1_IN 0
`define FSI4RXD1_OE 0
`define FSI4RXD1_OUT 0
`define FSI4TXCLK_IN 0
`define FSI4TXCLK_OE 0
`define FSI4TXCLK_OUT 0
`define FSI4TXD0_IN 0
`define FSI4TXD0_OE 0
`define FSI4TXD0_OUT 0
`define FSI4TXD1_IN 0
`define FSI4TXD1_OE 0
`define FSI4TXD1_OUT 0
`define FSI5RXCLK_IN 0
`define FSI5RXCLK_OE 0
`define FSI5RXCLK_OUT 0
`define FSI5RXD0_IN 0
`define FSI5RXD0_OE 0
`define FSI5RXD0_OUT 0
`define FSI5RXD1_IN 0
`define FSI5RXD1_OE 0
`define FSI5RXD1_OUT 0
`define FSI5TXCLK_IN 0
`define FSI5TXCLK_OE 0
`define FSI5TXCLK_OUT 0
`define FSI5TXD0_IN 0
`define FSI5TXD0_OE 0
`define FSI5TXD0_OUT 0
`define FSI5TXD1_IN 0
`define FSI5TXD1_OE 0
`define FSI5TXD1_OUT 0
`define GMII_MDC_IN 0
`define GMII_MDC_OE 0
`define GMII_MDC_OUT 0
`define GMII_MDIO_IN 0
`define GMII_MDIO_OE 0
`define GMII_MDIO_OUT 0
`define I2C0SCL_IN 0
`define I2C0SCL_OE 0
`define I2C0SCL_OUT 0
`define I2C0SDA_IN 0
`define I2C0SDA_OE 0
`define I2C0SDA_OUT 0
`define I2C1SCL_IN 0
`define I2C1SCL_OE 0
`define I2C1SCL_OUT 0
`define I2C1SDA_IN 0
`define I2C1SDA_OE 0
`define I2C1SDA_OUT 0
`define I2C2SCL_IN 0
`define I2C2SCL_OE 0
`define I2C2SCL_OUT 0
`define I2C2SDA_IN 0
`define I2C2SDA_OE 0
`define I2C2SDA_OUT 0
`define I2C3SCL_IN 0
`define I2C3SCL_OE 0
`define I2C3SCL_OUT 0
`define I2C3SDA_IN 0
`define I2C3SDA_OE 0
`define I2C3SDA_OUT 0
`define LIN0RX_IN 0
`define LIN0RX_OE 0
`define LIN0RX_OUT 0
`define LIN0TX_IN 0
`define LIN0TX_OE 0
`define LIN0TX_OUT 0
`define LIN1RX_IN 0
`define LIN1RX_OE 0
`define LIN1RX_OUT 0
`define LIN1TX_IN 0
`define LIN1TX_OE 0
`define LIN1TX_OUT 0
`define LIN2RX_IN 0
`define LIN2RX_OE 0
`define LIN2RX_OUT 0
`define LIN2TX_IN 0
`define LIN2TX_OE 0
`define LIN2TX_OUT 0
`define LIN3RX_IN 0
`define LIN3RX_OE 0
`define LIN3RX_OUT 0
`define LIN3TX_IN 0
`define LIN3TX_OE 0
`define LIN3TX_OUT 0
`define LIN4RX_IN 0
`define LIN4RX_OE 0
`define LIN4RX_OUT 0
`define LIN4TX_IN 0
`define LIN4TX_OE 0
`define LIN4TX_OUT 0
`define LIN5RX_IN 0
`define LIN5RX_OE 0
`define LIN5RX_OUT 0
`define LIN5TX_IN 0
`define LIN5TX_OE 0
`define LIN5TX_OUT 0
`define LIN6RX_IN 0
`define LIN6RX_OE 0
`define LIN6RX_OUT 0
`define LIN6TX_IN 0
`define LIN6TX_OE 0
`define LIN6TX_OUT 0
`define LIN7RX_IN 0
`define LIN7RX_OE 0
`define LIN7RX_OUT 0
`define LIN7TX_IN 0
`define LIN7TX_OE 0
`define LIN7TX_OUT 0
`define LPD_A_PWM1A_IN 0
`define LPD_A_PWM1A_OE 0
`define LPD_A_PWM1A_OUT 0
`define LPD_A_PWM1B_IN 0
`define LPD_A_PWM1B_OE 0
`define LPD_A_PWM1B_OUT 0
`define LPD_A_PWM2A_IN 0
`define LPD_A_PWM2A_OE 0
`define LPD_A_PWM2A_OUT 0
`define LPD_A_PWM2B_IN 0
`define LPD_A_PWM2B_OE 0
`define LPD_A_PWM2B_OUT 0
`define LPD_B_PWM3A_IN 0
`define LPD_B_PWM3A_OE 0
`define LPD_B_PWM3A_OUT 0
`define LPD_B_PWM3B_IN 0
`define LPD_B_PWM3B_OE 0
`define LPD_B_PWM3B_OUT 0
`define LPD_B_PWM4A_IN 0
`define LPD_B_PWM4A_OE 0
`define LPD_B_PWM4A_OUT 0
`define LPD_B_PWM4B_IN 0
`define LPD_B_PWM4B_OE 0
`define LPD_B_PWM4B_OUT 0
`define LPD_CAN0RX_IN 0
`define LPD_CAN0RX_OE 0
`define LPD_CAN0RX_OUT 0
`define LPD_CAN0TX_IN 0
`define LPD_CAN0TX_OE 0
`define LPD_CAN0TX_OUT 0
`define LPD_LIN0RX_IN 0
`define LPD_LIN0RX_OE 0
`define LPD_LIN0RX_OUT 0
`define LPD_LIN0TX_IN 0
`define LPD_LIN0TX_OE 0
`define LPD_LIN0TX_OUT 0
`define MCASP0ACLKR_IN 0
`define MCASP0ACLKR_OE 0
`define MCASP0ACLKR_OUT 0
`define MCASP0ACLKX_IN 0
`define MCASP0ACLKX_OE 0
`define MCASP0ACLKX_OUT 0
`define MCASP0AFSR_IN 0
`define MCASP0AFSR_OE 0
`define MCASP0AFSR_OUT 0
`define MCASP0AFSX_IN 0
`define MCASP0AFSX_OE 0
`define MCASP0AFSX_OUT 0
`define MCASP0AXR0_IN 0
`define MCASP0AXR0_OE 0
`define MCASP0AXR0_OUT 0
`define MCASP0AXR1_IN 0
`define MCASP0AXR1_OE 0
`define MCASP0AXR1_OUT 0
`define MCASP0AXR2_IN 0
`define MCASP0AXR2_OE 0
`define MCASP0AXR2_OUT 0
`define MCASP0AXR3_IN 0
`define MCASP0AXR3_OE 0
`define MCASP0AXR3_OUT 0
`define MCASP0EXTREFCLK_IN 0
`define MCASP0EXTREFCLK_OE 0
`define MCASP0EXTREFCLK_OUT 0
`define MCPWM0A_IN 0
`define MCPWM0A_OE 0
`define MCPWM0A_OUT 0
`define MCPWM0B_IN 0
`define MCPWM0B_OE 0
`define MCPWM0B_OUT 0
`define MCPWM0C_IN 0
`define MCPWM0C_OE 0
`define MCPWM0C_OUT 0
`define MCPWM0D_IN 0
`define MCPWM0D_OE 0
`define MCPWM0D_OUT 0
`define MCPWM0E_IN 0
`define MCPWM0E_OE 0
`define MCPWM0E_OUT 0
`define MCPWM0F_IN 0
`define MCPWM0F_OE 0
`define MCPWM0F_OUT 0
`define MCPWM10A_IN 0
`define MCPWM10A_OE 0
`define MCPWM10A_OUT 0
`define MCPWM10B_IN 0
`define MCPWM10B_OE 0
`define MCPWM10B_OUT 0
`define MCPWM10C_IN 0
`define MCPWM10C_OE 0
`define MCPWM10C_OUT 0
`define MCPWM10D_IN 0
`define MCPWM10D_OE 0
`define MCPWM10D_OUT 0
`define MCPWM10E_IN 0
`define MCPWM10E_OE 0
`define MCPWM10E_OUT 0
`define MCPWM10F_IN 0
`define MCPWM10F_OE 0
`define MCPWM10F_OUT 0
`define MCPWM1A_IN 0
`define MCPWM1A_OE 0
`define MCPWM1A_OUT 0
`define MCPWM1B_IN 0
`define MCPWM1B_OE 0
`define MCPWM1B_OUT 0
`define MCPWM1C_IN 0
`define MCPWM1C_OE 0
`define MCPWM1C_OUT 0
`define MCPWM1D_IN 0
`define MCPWM1D_OE 0
`define MCPWM1D_OUT 0
`define MCPWM1E_IN 0
`define MCPWM1E_OE 0
`define MCPWM1E_OUT 0
`define MCPWM1F_IN 0
`define MCPWM1F_OE 0
`define MCPWM1F_OUT 0
`define MCPWM2A_IN 0
`define MCPWM2A_OE 0
`define MCPWM2A_OUT 0
`define MCPWM2B_IN 0
`define MCPWM2B_OE 0
`define MCPWM2B_OUT 0
`define MCPWM2C_IN 0
`define MCPWM2C_OE 0
`define MCPWM2C_OUT 0
`define MCPWM2D_IN 0
`define MCPWM2D_OE 0
`define MCPWM2D_OUT 0
`define MCPWM2E_IN 0
`define MCPWM2E_OE 0
`define MCPWM2E_OUT 0
`define MCPWM2F_IN 0
`define MCPWM2F_OE 0
`define MCPWM2F_OUT 0
`define MCPWM3A_IN 0
`define MCPWM3A_OE 0
`define MCPWM3A_OUT 0
`define MCPWM3B_IN 0
`define MCPWM3B_OE 0
`define MCPWM3B_OUT 0
`define MCPWM3C_IN 0
`define MCPWM3C_OE 0
`define MCPWM3C_OUT 0
`define MCPWM3D_IN 0
`define MCPWM3D_OE 0
`define MCPWM3D_OUT 0
`define MCPWM3E_IN 0
`define MCPWM3E_OE 0
`define MCPWM3E_OUT 0
`define MCPWM3F_IN 0
`define MCPWM3F_OE 0
`define MCPWM3F_OUT 0
`define MCPWM4A_IN 0
`define MCPWM4A_OE 0
`define MCPWM4A_OUT 0
`define MCPWM4B_IN 0
`define MCPWM4B_OE 0
`define MCPWM4B_OUT 0
`define MCPWM4C_IN 0
`define MCPWM4C_OE 0
`define MCPWM4C_OUT 0
`define MCPWM4D_IN 0
`define MCPWM4D_OE 0
`define MCPWM4D_OUT 0
`define MCPWM4E_IN 0
`define MCPWM4E_OE 0
`define MCPWM4E_OUT 0
`define MCPWM4F_IN 0
`define MCPWM4F_OE 0
`define MCPWM4F_OUT 0
`define MCPWM5A_IN 0
`define MCPWM5A_OE 0
`define MCPWM5A_OUT 0
`define MCPWM5B_IN 0
`define MCPWM5B_OE 0
`define MCPWM5B_OUT 0
`define MCPWM5C_IN 0
`define MCPWM5C_OE 0
`define MCPWM5C_OUT 0
`define MCPWM5D_IN 0
`define MCPWM5D_OE 0
`define MCPWM5D_OUT 0
`define MCPWM5E_IN 0
`define MCPWM5E_OE 0
`define MCPWM5E_OUT 0
`define MCPWM5F_IN 0
`define MCPWM5F_OE 0
`define MCPWM5F_OUT 0
`define MCPWM6A_IN 0
`define MCPWM6A_OE 0
`define MCPWM6A_OUT 0
`define MCPWM6B_IN 0
`define MCPWM6B_OE 0
`define MCPWM6B_OUT 0
`define MCPWM6C_IN 0
`define MCPWM6C_OE 0
`define MCPWM6C_OUT 0
`define MCPWM6D_IN 0
`define MCPWM6D_OE 0
`define MCPWM6D_OUT 0
`define MCPWM6E_IN 0
`define MCPWM6E_OE 0
`define MCPWM6E_OUT 0
`define MCPWM6F_IN 0
`define MCPWM6F_OE 0
`define MCPWM6F_OUT 0
`define MCPWM7A_IN 0
`define MCPWM7A_OE 0
`define MCPWM7A_OUT 0
`define MCPWM7B_IN 0
`define MCPWM7B_OE 0
`define MCPWM7B_OUT 0
`define MCPWM7C_IN 0
`define MCPWM7C_OE 0
`define MCPWM7C_OUT 0
`define MCPWM7D_IN 0
`define MCPWM7D_OE 0
`define MCPWM7D_OUT 0
`define MCPWM7E_IN 0
`define MCPWM7E_OE 0
`define MCPWM7E_OUT 0
`define MCPWM7F_IN 0
`define MCPWM7F_OE 0
`define MCPWM7F_OUT 0
`define MCPWM8A_IN 0
`define MCPWM8A_OE 0
`define MCPWM8A_OUT 0
`define MCPWM8B_IN 0
`define MCPWM8B_OE 0
`define MCPWM8B_OUT 0
`define MCPWM8C_IN 0
`define MCPWM8C_OE 0
`define MCPWM8C_OUT 0
`define MCPWM8D_IN 0
`define MCPWM8D_OE 0
`define MCPWM8D_OUT 0
`define MCPWM8E_IN 0
`define MCPWM8E_OE 0
`define MCPWM8E_OUT 0
`define MCPWM8F_IN 0
`define MCPWM8F_OE 0
`define MCPWM8F_OUT 0
`define MCPWM9A_IN 0
`define MCPWM9A_OE 0
`define MCPWM9A_OUT 0
`define MCPWM9B_IN 0
`define MCPWM9B_OE 0
`define MCPWM9B_OUT 0
`define MCPWM9C_IN 0
`define MCPWM9C_OE 0
`define MCPWM9C_OUT 0
`define MCPWM9D_IN 0
`define MCPWM9D_OE 0
`define MCPWM9D_OUT 0
`define MCPWM9E_IN 0
`define MCPWM9E_OE 0
`define MCPWM9E_OUT 0
`define MCPWM9F_IN 0
`define MCPWM9F_OE 0
`define MCPWM9F_OUT 0
`define MIBSPI0CLK_IN 0
`define MIBSPI0CLK_OE 0
`define MIBSPI0CLK_OUT 0
`define MIBSPI0CS0_IN 0
`define MIBSPI0CS0_OE 0
`define MIBSPI0CS0_OUT 0
`define MIBSPI0CS10_IN 0
`define MIBSPI0CS10_OE 0
`define MIBSPI0CS10_OUT 0
`define MIBSPI0CS11_IN 0
`define MIBSPI0CS11_OE 0
`define MIBSPI0CS11_OUT 0
`define MIBSPI0CS1_IN 0
`define MIBSPI0CS1_OE 0
`define MIBSPI0CS1_OUT 0
`define MIBSPI0CS2_IN 0
`define MIBSPI0CS2_OE 0
`define MIBSPI0CS2_OUT 0
`define MIBSPI0CS3_IN 0
`define MIBSPI0CS3_OE 0
`define MIBSPI0CS3_OUT 0
`define MIBSPI0CS4_IN 0
`define MIBSPI0CS4_OE 0
`define MIBSPI0CS4_OUT 0
`define MIBSPI0CS5_IN 0
`define MIBSPI0CS5_OE 0
`define MIBSPI0CS5_OUT 0
`define MIBSPI0CS6_IN 0
`define MIBSPI0CS6_OE 0
`define MIBSPI0CS6_OUT 0
`define MIBSPI0CS7_IN 0
`define MIBSPI0CS7_OE 0
`define MIBSPI0CS7_OUT 0
`define MIBSPI0CS8_IN 0
`define MIBSPI0CS8_OE 0
`define MIBSPI0CS8_OUT 0
`define MIBSPI0CS9_IN 0
`define MIBSPI0CS9_OE 0
`define MIBSPI0CS9_OUT 0
`define MIBSPI0PICO_IN 0
`define MIBSPI0PICO_OE 0
`define MIBSPI0PICO_OUT 0
`define MIBSPI0POCI_IN 0
`define MIBSPI0POCI_OE 0
`define MIBSPI0POCI_OUT 0
`define MIBSPI1CLK_IN 0
`define MIBSPI1CLK_OE 0
`define MIBSPI1CLK_OUT 0
`define MIBSPI1CS0_IN 0
`define MIBSPI1CS0_OE 0
`define MIBSPI1CS0_OUT 0
`define MIBSPI1CS10_IN 0
`define MIBSPI1CS10_OE 0
`define MIBSPI1CS10_OUT 0
`define MIBSPI1CS11_IN 0
`define MIBSPI1CS11_OE 0
`define MIBSPI1CS11_OUT 0
`define MIBSPI1CS1_IN 0
`define MIBSPI1CS1_OE 0
`define MIBSPI1CS1_OUT 0
`define MIBSPI1CS2_IN 0
`define MIBSPI1CS2_OE 0
`define MIBSPI1CS2_OUT 0
`define MIBSPI1CS3_IN 0
`define MIBSPI1CS3_OE 0
`define MIBSPI1CS3_OUT 0
`define MIBSPI1CS4_IN 0
`define MIBSPI1CS4_OE 0
`define MIBSPI1CS4_OUT 0
`define MIBSPI1CS5_IN 0
`define MIBSPI1CS5_OE 0
`define MIBSPI1CS5_OUT 0
`define MIBSPI1CS6_IN 0
`define MIBSPI1CS6_OE 0
`define MIBSPI1CS6_OUT 0
`define MIBSPI1CS7_IN 0
`define MIBSPI1CS7_OE 0
`define MIBSPI1CS7_OUT 0
`define MIBSPI1CS8_IN 0
`define MIBSPI1CS8_OE 0
`define MIBSPI1CS8_OUT 0
`define MIBSPI1CS9_IN 0
`define MIBSPI1CS9_OE 0
`define MIBSPI1CS9_OUT 0
`define MIBSPI1PICO_IN 0
`define MIBSPI1PICO_OE 0
`define MIBSPI1PICO_OUT 0
`define MIBSPI1POCI_IN 0
`define MIBSPI1POCI_OE 0
`define MIBSPI1POCI_OUT 0
`define MMC0CD_IN 0
`define MMC0CD_OE 0
`define MMC0CD_OUT 0
`define MMC0CLK_IN 0
`define MMC0CLK_OE 0
`define MMC0CLK_OUT 0
`define MMC0CMD_IN 0
`define MMC0CMD_OE 0
`define MMC0CMD_OUT 0
`define MMC0DATA0_IN 0
`define MMC0DATA0_OE 0
`define MMC0DATA0_OUT 0
`define MMC0DATA1_IN 0
`define MMC0DATA1_OE 0
`define MMC0DATA1_OUT 0
`define MMC0DATA2_IN 0
`define MMC0DATA2_OE 0
`define MMC0DATA2_OUT 0
`define MMC0DATA3_IN 0
`define MMC0DATA3_OE 0
`define MMC0DATA3_OUT 0
`define MMC0WP_IN 0
`define MMC0WP_OE 0
`define MMC0WP_OUT 0
`define MP0_0 0
`define MP0_0_GPIO_OUTPUT_ENABLE 0
`define MP0_0_INFUNC_EN 0
`define MP0_0_OUTFUNC_SEL 0
`define MP0_0_PINCTRL_0_IE 0
`define MP0_0_PINCTRL_0_OD 0
`define MP0_0_PULLEN 0
`define MP0_0_PULLSEL 0
`define MP0_0_pad_y 0
`define MP0_1 0
`define MP0_10 0
`define MP0_10_GPIO_OUTPUT_ENABLE 0
`define MP0_10_INFUNC_EN 0
`define MP0_10_OUTFUNC_SEL 0
`define MP0_10_PINCTRL_0_IE 0
`define MP0_10_PINCTRL_0_OD 0
`define MP0_10_PULLEN 0
`define MP0_10_PULLSEL 0
`define MP0_10_pad_y 0
`define MP0_11 0
`define MP0_11_GPIO_OUTPUT_ENABLE 0
`define MP0_11_INFUNC_EN 0
`define MP0_11_OUTFUNC_SEL 0
`define MP0_11_PINCTRL_0_IE 0
`define MP0_11_PINCTRL_0_OD 0
`define MP0_11_PULLEN 0
`define MP0_11_PULLSEL 0
`define MP0_11_pad_y 0
`define MP0_12 0
`define MP0_12_GPIO_OUTPUT_ENABLE 0
`define MP0_12_INFUNC_EN 0
`define MP0_12_OUTFUNC_SEL 0
`define MP0_12_PINCTRL_0_IE 0
`define MP0_12_PINCTRL_0_OD 0
`define MP0_12_PULLEN 0
`define MP0_12_PULLSEL 0
`define MP0_12_pad_y 0
`define MP0_13 0
`define MP0_13_GPIO_OUTPUT_ENABLE 0
`define MP0_13_INFUNC_EN 0
`define MP0_13_OUTFUNC_SEL 0
`define MP0_13_PINCTRL_0_IE 0
`define MP0_13_PINCTRL_0_OD 0
`define MP0_13_PULLEN 0
`define MP0_13_PULLSEL 0
`define MP0_13_pad_y 0
`define MP0_14 0
`define MP0_14_GPIO_OUTPUT_ENABLE 0
`define MP0_14_INFUNC_EN 0
`define MP0_14_OUTFUNC_SEL 0
`define MP0_14_PINCTRL_0_IE 0
`define MP0_14_PINCTRL_0_OD 0
`define MP0_14_PULLEN 0
`define MP0_14_PULLSEL 0
`define MP0_14_pad_y 0
`define MP0_15 0
`define MP0_15_GPIO_OUTPUT_ENABLE 0
`define MP0_15_INFUNC_EN 0
`define MP0_15_OUTFUNC_SEL 0
`define MP0_15_PINCTRL_0_IE 0
`define MP0_15_PINCTRL_0_OD 0
`define MP0_15_PULLEN 0
`define MP0_15_PULLSEL 0
`define MP0_15_pad_y 0
`define MP0_16 0
`define MP0_16_GPIO_OUTPUT_ENABLE 0
`define MP0_16_INFUNC_EN 0
`define MP0_16_OUTFUNC_SEL 0
`define MP0_16_PINCTRL_0_IE 0
`define MP0_16_PINCTRL_0_OD 0
`define MP0_16_PULLEN 0
`define MP0_16_PULLSEL 0
`define MP0_16_pad_y 0
`define MP0_17 0
`define MP0_17_GPIO_OUTPUT_ENABLE 0
`define MP0_17_INFUNC_EN 0
`define MP0_17_OUTFUNC_SEL 0
`define MP0_17_PINCTRL_0_IE 0
`define MP0_17_PINCTRL_0_OD 0
`define MP0_17_PULLEN 0
`define MP0_17_PULLSEL 0
`define MP0_17_pad_y 0
`define MP0_18 0
`define MP0_18_GPIO_OUTPUT_ENABLE 0
`define MP0_18_INFUNC_EN 0
`define MP0_18_OUTFUNC_SEL 0
`define MP0_18_PINCTRL_0_IE 0
`define MP0_18_PINCTRL_0_OD 0
`define MP0_18_PULLEN 0
`define MP0_18_PULLSEL 0
`define MP0_18_pad_y 0
`define MP0_19 0
`define MP0_19_GPIO_OUTPUT_ENABLE 0
`define MP0_19_INFUNC_EN 0
`define MP0_19_OUTFUNC_SEL 0
`define MP0_19_PINCTRL_0_IE 0
`define MP0_19_PINCTRL_0_OD 0
`define MP0_19_PULLEN 0
`define MP0_19_PULLSEL 0
`define MP0_19_pad_y 0
`define MP0_1_GPIO_OUTPUT_ENABLE 0
`define MP0_1_INFUNC_EN 0
`define MP0_1_OUTFUNC_SEL 0
`define MP0_1_PINCTRL_0_IE 0
`define MP0_1_PINCTRL_0_OD 0
`define MP0_1_PULLEN 0
`define MP0_1_PULLSEL 0
`define MP0_1_pad_y 0
`define MP0_2 0
`define MP0_20 0
`define MP0_20_GPIO_OUTPUT_ENABLE 0
`define MP0_20_INFUNC_EN 0
`define MP0_20_OUTFUNC_SEL 0
`define MP0_20_PINCTRL_0_IE 0
`define MP0_20_PINCTRL_0_OD 0
`define MP0_20_PULLEN 0
`define MP0_20_PULLSEL 0
`define MP0_20_pad_y 0
`define MP0_21 0
`define MP0_21_GPIO_OUTPUT_ENABLE 0
`define MP0_21_INFUNC_EN 0
`define MP0_21_OUTFUNC_SEL 0
`define MP0_21_PINCTRL_0_IE 0
`define MP0_21_PINCTRL_0_OD 0
`define MP0_21_PULLEN 0
`define MP0_21_PULLSEL 0
`define MP0_21_pad_y 0
`define MP0_22 0
`define MP0_22_GPIO_OUTPUT_ENABLE 0
`define MP0_22_INFUNC_EN 0
`define MP0_22_OUTFUNC_SEL 0
`define MP0_22_PINCTRL_0_IE 0
`define MP0_22_PINCTRL_0_OD 0
`define MP0_22_PULLEN 0
`define MP0_22_PULLSEL 0
`define MP0_22_pad_y 0
`define MP0_23 0
`define MP0_23_GPIO_OUTPUT_ENABLE 0
`define MP0_23_INFUNC_EN 0
`define MP0_23_OUTFUNC_SEL 0
`define MP0_23_PINCTRL_0_IE 0
`define MP0_23_PINCTRL_0_OD 0
`define MP0_23_PULLEN 0
`define MP0_23_PULLSEL 0
`define MP0_23_pad_y 0
`define MP0_24 0
`define MP0_24_GPIO_OUTPUT_ENABLE 0
`define MP0_24_INFUNC_EN 0
`define MP0_24_OUTFUNC_SEL 0
`define MP0_24_PINCTRL_0_IE 0
`define MP0_24_PINCTRL_0_OD 0
`define MP0_24_PULLEN 0
`define MP0_24_PULLSEL 0
`define MP0_24_pad_y 0
`define MP0_25 0
`define MP0_25_GPIO_OUTPUT_ENABLE 0
`define MP0_25_INFUNC_EN 0
`define MP0_25_OUTFUNC_SEL 0
`define MP0_25_PINCTRL_0_IE 0
`define MP0_25_PINCTRL_0_OD 0
`define MP0_25_PULLEN 0
`define MP0_25_PULLSEL 0
`define MP0_25_pad_y 0
`define MP0_26 0
`define MP0_26_GPIO_OUTPUT_ENABLE 0
`define MP0_26_INFUNC_EN 0
`define MP0_26_OUTFUNC_SEL 0
`define MP0_26_PINCTRL_0_IE 0
`define MP0_26_PINCTRL_0_OD 0
`define MP0_26_PULLEN 0
`define MP0_26_PULLSEL 0
`define MP0_26_pad_y 0
`define MP0_27 0
`define MP0_27_GPIO_OUTPUT_ENABLE 0
`define MP0_27_INFUNC_EN 0
`define MP0_27_OUTFUNC_SEL 0
`define MP0_27_PINCTRL_0_IE 0
`define MP0_27_PINCTRL_0_OD 0
`define MP0_27_PULLEN 0
`define MP0_27_PULLSEL 0
`define MP0_27_pad_y 0
`define MP0_28 0
`define MP0_28_GPIO_OUTPUT_ENABLE 0
`define MP0_28_INFUNC_EN 0
`define MP0_28_OUTFUNC_SEL 0
`define MP0_28_PINCTRL_0_IE 0
`define MP0_28_PINCTRL_0_OD 0
`define MP0_28_PULLEN 0
`define MP0_28_PULLSEL 0
`define MP0_28_pad_y 0
`define MP0_29 0
`define MP0_29_GPIO_OUTPUT_ENABLE 0
`define MP0_29_INFUNC_EN 0
`define MP0_29_OUTFUNC_SEL 0
`define MP0_29_PINCTRL_0_IE 0
`define MP0_29_PINCTRL_0_OD 0
`define MP0_29_PULLEN 0
`define MP0_29_PULLSEL 0
`define MP0_29_pad_y 0
`define MP0_2_GPIO_OUTPUT_ENABLE 0
`define MP0_2_INFUNC_EN 0
`define MP0_2_OUTFUNC_SEL 0
`define MP0_2_PINCTRL_0_IE 0
`define MP0_2_PINCTRL_0_OD 0
`define MP0_2_PULLEN 0
`define MP0_2_PULLSEL 0
`define MP0_2_pad_y 0
`define MP0_3 0
`define MP0_30 0
`define MP0_30_GPIO_OUTPUT_ENABLE 0
`define MP0_30_INFUNC_EN 0
`define MP0_30_OUTFUNC_SEL 0
`define MP0_30_PINCTRL_0_IE 0
`define MP0_30_PINCTRL_0_OD 0
`define MP0_30_PULLEN 0
`define MP0_30_PULLSEL 0
`define MP0_30_pad_y 0
`define MP0_31 0
`define MP0_31_GPIO_OUTPUT_ENABLE 0
`define MP0_31_INFUNC_EN 0
`define MP0_31_OUTFUNC_SEL 0
`define MP0_31_PINCTRL_0_IE 0
`define MP0_31_PINCTRL_0_OD 0
`define MP0_31_PULLEN 0
`define MP0_31_PULLSEL 0
`define MP0_31_pad_y 0
`define MP0_3_GPIO_OUTPUT_ENABLE 0
`define MP0_3_INFUNC_EN 0
`define MP0_3_OUTFUNC_SEL 0
`define MP0_3_PINCTRL_0_IE 0
`define MP0_3_PINCTRL_0_OD 0
`define MP0_3_PULLEN 0
`define MP0_3_PULLSEL 0
`define MP0_3_pad_y 0
`define MP0_4 0
`define MP0_4_GPIO_OUTPUT_ENABLE 0
`define MP0_4_INFUNC_EN 0
`define MP0_4_OUTFUNC_SEL 0
`define MP0_4_PINCTRL_0_IE 0
`define MP0_4_PINCTRL_0_OD 0
`define MP0_4_PULLEN 0
`define MP0_4_PULLSEL 0
`define MP0_4_pad_y 0
`define MP0_5 0
`define MP0_5_GPIO_OUTPUT_ENABLE 0
`define MP0_5_INFUNC_EN 0
`define MP0_5_OUTFUNC_SEL 0
`define MP0_5_PINCTRL_0_IE 0
`define MP0_5_PINCTRL_0_OD 0
`define MP0_5_PULLEN 0
`define MP0_5_PULLSEL 0
`define MP0_5_pad_y 0
`define MP0_6 0
`define MP0_6_GPIO_OUTPUT_ENABLE 0
`define MP0_6_INFUNC_EN 0
`define MP0_6_OUTFUNC_SEL 0
`define MP0_6_PINCTRL_0_IE 0
`define MP0_6_PINCTRL_0_OD 0
`define MP0_6_PULLEN 0
`define MP0_6_PULLSEL 0
`define MP0_6_pad_y 0
`define MP0_7 0
`define MP0_7_GPIO_OUTPUT_ENABLE 0
`define MP0_7_INFUNC_EN 0
`define MP0_7_OUTFUNC_SEL 0
`define MP0_7_PINCTRL_0_IE 0
`define MP0_7_PINCTRL_0_OD 0
`define MP0_7_PULLEN 0
`define MP0_7_PULLSEL 0
`define MP0_7_pad_y 0
`define MP0_8 0
`define MP0_8_GPIO_OUTPUT_ENABLE 0
`define MP0_8_INFUNC_EN 0
`define MP0_8_OUTFUNC_SEL 0
`define MP0_8_PINCTRL_0_IE 0
`define MP0_8_PINCTRL_0_OD 0
`define MP0_8_PULLEN 0
`define MP0_8_PULLSEL 0
`define MP0_8_pad_y 0
`define MP0_9 0
`define MP0_9_GPIO_OUTPUT_ENABLE 0
`define MP0_9_INFUNC_EN 0
`define MP0_9_OUTFUNC_SEL 0
`define MP0_9_PINCTRL_0_IE 0
`define MP0_9_PINCTRL_0_OD 0
`define MP0_9_PULLEN 0
`define MP0_9_PULLSEL 0
`define MP0_9_pad_y 0
`define MP1_0 0
`define MP1_0_GPIO_OUTPUT_ENABLE 0
`define MP1_0_INFUNC_EN 0
`define MP1_0_OUTFUNC_SEL 0
`define MP1_0_PINCTRL_0_IE 0
`define MP1_0_PINCTRL_0_OD 0
`define MP1_0_PULLEN 0
`define MP1_0_PULLSEL 0
`define MP1_0_pad_y 0
`define MP1_1 0
`define MP1_10 0
`define MP1_10_GPIO_OUTPUT_ENABLE 0
`define MP1_10_INFUNC_EN 0
`define MP1_10_OUTFUNC_SEL 0
`define MP1_10_PINCTRL_0_IE 0
`define MP1_10_PINCTRL_0_OD 0
`define MP1_10_PULLEN 0
`define MP1_10_PULLSEL 0
`define MP1_10_pad_y 0
`define MP1_11 0
`define MP1_11_GPIO_OUTPUT_ENABLE 0
`define MP1_11_INFUNC_EN 0
`define MP1_11_OUTFUNC_SEL 0
`define MP1_11_PINCTRL_0_IE 0
`define MP1_11_PINCTRL_0_OD 0
`define MP1_11_PULLEN 0
`define MP1_11_PULLSEL 0
`define MP1_11_pad_y 0
`define MP1_12 0
`define MP1_12_GPIO_OUTPUT_ENABLE 0
`define MP1_12_INFUNC_EN 0
`define MP1_12_OUTFUNC_SEL 0
`define MP1_12_PINCTRL_0_IE 0
`define MP1_12_PINCTRL_0_OD 0
`define MP1_12_PULLEN 0
`define MP1_12_PULLSEL 0
`define MP1_12_pad_y 0
`define MP1_13 0
`define MP1_13_GPIO_OUTPUT_ENABLE 0
`define MP1_13_INFUNC_EN 0
`define MP1_13_OUTFUNC_SEL 0
`define MP1_13_PINCTRL_0_IE 0
`define MP1_13_PINCTRL_0_OD 0
`define MP1_13_PULLEN 0
`define MP1_13_PULLSEL 0
`define MP1_13_pad_y 0
`define MP1_14 0
`define MP1_14_GPIO_OUTPUT_ENABLE 0
`define MP1_14_INFUNC_EN 0
`define MP1_14_OUTFUNC_SEL 0
`define MP1_14_PINCTRL_0_IE 0
`define MP1_14_PINCTRL_0_OD 0
`define MP1_14_PULLEN 0
`define MP1_14_PULLSEL 0
`define MP1_14_pad_y 0
`define MP1_15 0
`define MP1_15_GPIO_OUTPUT_ENABLE 0
`define MP1_15_INFUNC_EN 0
`define MP1_15_OUTFUNC_SEL 0
`define MP1_15_PINCTRL_0_IE 0
`define MP1_15_PINCTRL_0_OD 0
`define MP1_15_PULLEN 0
`define MP1_15_PULLSEL 0
`define MP1_15_pad_y 0
`define MP1_1_GPIO_OUTPUT_ENABLE 0
`define MP1_1_INFUNC_EN 0
`define MP1_1_OUTFUNC_SEL 0
`define MP1_1_PINCTRL_0_IE 0
`define MP1_1_PINCTRL_0_OD 0
`define MP1_1_PULLEN 0
`define MP1_1_PULLSEL 0
`define MP1_1_pad_y 0
`define MP1_2 0
`define MP1_2_GPIO_OUTPUT_ENABLE 0
`define MP1_2_INFUNC_EN 0
`define MP1_2_OUTFUNC_SEL 0
`define MP1_2_PINCTRL_0_IE 0
`define MP1_2_PINCTRL_0_OD 0
`define MP1_2_PULLEN 0
`define MP1_2_PULLSEL 0
`define MP1_2_pad_y 0
`define MP1_3 0
`define MP1_3_GPIO_OUTPUT_ENABLE 0
`define MP1_3_INFUNC_EN 0
`define MP1_3_OUTFUNC_SEL 0
`define MP1_3_PINCTRL_0_IE 0
`define MP1_3_PINCTRL_0_OD 0
`define MP1_3_PULLEN 0
`define MP1_3_PULLSEL 0
`define MP1_3_pad_y 0
`define MP1_4 0
`define MP1_4_GPIO_OUTPUT_ENABLE 0
`define MP1_4_INFUNC_EN 0
`define MP1_4_OUTFUNC_SEL 0
`define MP1_4_PINCTRL_0_IE 0
`define MP1_4_PINCTRL_0_OD 0
`define MP1_4_PULLEN 0
`define MP1_4_PULLSEL 0
`define MP1_4_pad_y 0
`define MP1_5 0
`define MP1_5_GPIO_OUTPUT_ENABLE 0
`define MP1_5_INFUNC_EN 0
`define MP1_5_OUTFUNC_SEL 0
`define MP1_5_PINCTRL_0_IE 0
`define MP1_5_PINCTRL_0_OD 0
`define MP1_5_PULLEN 0
`define MP1_5_PULLSEL 0
`define MP1_5_pad_y 0
`define MP1_6 0
`define MP1_6_GPIO_OUTPUT_ENABLE 0
`define MP1_6_INFUNC_EN 0
`define MP1_6_OUTFUNC_SEL 0
`define MP1_6_PINCTRL_0_IE 0
`define MP1_6_PINCTRL_0_OD 0
`define MP1_6_PULLEN 0
`define MP1_6_PULLSEL 0
`define MP1_6_pad_y 0
`define MP1_7 0
`define MP1_7_GPIO_OUTPUT_ENABLE 0
`define MP1_7_INFUNC_EN 0
`define MP1_7_OUTFUNC_SEL 0
`define MP1_7_PINCTRL_0_IE 0
`define MP1_7_PINCTRL_0_OD 0
`define MP1_7_PULLEN 0
`define MP1_7_PULLSEL 0
`define MP1_7_pad_y 0
`define MP1_8 0
`define MP1_8_GPIO_OUTPUT_ENABLE 0
`define MP1_8_INFUNC_EN 0
`define MP1_8_OUTFUNC_SEL 0
`define MP1_8_PINCTRL_0_IE 0
`define MP1_8_PINCTRL_0_OD 0
`define MP1_8_PULLEN 0
`define MP1_8_PULLSEL 0
`define MP1_8_pad_y 0
`define MP1_9 0
`define MP1_9_GPIO_OUTPUT_ENABLE 0
`define MP1_9_INFUNC_EN 0
`define MP1_9_OUTFUNC_SEL 0
`define MP1_9_PINCTRL_0_IE 0
`define MP1_9_PINCTRL_0_OD 0
`define MP1_9_PULLEN 0
`define MP1_9_PULLSEL 0
`define MP1_9_pad_y 0
`define MP2_0 0
`define MP2_0_GPIO_OUTPUT_ENABLE 0
`define MP2_0_INFUNC_EN 0
`define MP2_0_OUTFUNC_SEL 0
`define MP2_0_PINCTRL_0_IE 0
`define MP2_0_PINCTRL_0_OD 0
`define MP2_0_PULLEN 0
`define MP2_0_PULLSEL 0
`define MP2_0_pad_y 0
`define MP2_1 0
`define MP2_10 0
`define MP2_10_GPIO_OUTPUT_ENABLE 0
`define MP2_10_INFUNC_EN 0
`define MP2_10_OUTFUNC_SEL 0
`define MP2_10_PINCTRL_0_IE 0
`define MP2_10_PINCTRL_0_OD 0
`define MP2_10_PULLEN 0
`define MP2_10_PULLSEL 0
`define MP2_10_pad_y 0
`define MP2_11 0
`define MP2_11_GPIO_OUTPUT_ENABLE 0
`define MP2_11_INFUNC_EN 0
`define MP2_11_OUTFUNC_SEL 0
`define MP2_11_PINCTRL_0_IE 0
`define MP2_11_PINCTRL_0_OD 0
`define MP2_11_PULLEN 0
`define MP2_11_PULLSEL 0
`define MP2_11_pad_y 0
`define MP2_12 0
`define MP2_12_GPIO_OUTPUT_ENABLE 0
`define MP2_12_INFUNC_EN 0
`define MP2_12_OUTFUNC_SEL 0
`define MP2_12_PINCTRL_0_IE 0
`define MP2_12_PINCTRL_0_OD 0
`define MP2_12_PULLEN 0
`define MP2_12_PULLSEL 0
`define MP2_12_pad_y 0
`define MP2_13 0
`define MP2_13_GPIO_OUTPUT_ENABLE 0
`define MP2_13_INFUNC_EN 0
`define MP2_13_OUTFUNC_SEL 0
`define MP2_13_PINCTRL_0_IE 0
`define MP2_13_PINCTRL_0_OD 0
`define MP2_13_PULLEN 0
`define MP2_13_PULLSEL 0
`define MP2_13_pad_y 0
`define MP2_14 0
`define MP2_14_GPIO_OUTPUT_ENABLE 0
`define MP2_14_INFUNC_EN 0
`define MP2_14_OUTFUNC_SEL 0
`define MP2_14_PINCTRL_0_IE 0
`define MP2_14_PINCTRL_0_OD 0
`define MP2_14_PULLEN 0
`define MP2_14_PULLSEL 0
`define MP2_14_pad_y 0
`define MP2_15 0
`define MP2_15_GPIO_OUTPUT_ENABLE 0
`define MP2_15_INFUNC_EN 0
`define MP2_15_OUTFUNC_SEL 0
`define MP2_15_PINCTRL_0_IE 0
`define MP2_15_PINCTRL_0_OD 0
`define MP2_15_PULLEN 0
`define MP2_15_PULLSEL 0
`define MP2_15_pad_y 0
`define MP2_1_GPIO_OUTPUT_ENABLE 0
`define MP2_1_INFUNC_EN 0
`define MP2_1_OUTFUNC_SEL 0
`define MP2_1_PINCTRL_0_IE 0
`define MP2_1_PINCTRL_0_OD 0
`define MP2_1_PULLEN 0
`define MP2_1_PULLSEL 0
`define MP2_1_pad_y 0
`define MP2_2 0
`define MP2_2_GPIO_OUTPUT_ENABLE 0
`define MP2_2_INFUNC_EN 0
`define MP2_2_OUTFUNC_SEL 0
`define MP2_2_PINCTRL_0_IE 0
`define MP2_2_PINCTRL_0_OD 0
`define MP2_2_PULLEN 0
`define MP2_2_PULLSEL 0
`define MP2_2_pad_y 0
`define MP2_3 0
`define MP2_3_GPIO_OUTPUT_ENABLE 0
`define MP2_3_INFUNC_EN 0
`define MP2_3_OUTFUNC_SEL 0
`define MP2_3_PINCTRL_0_IE 0
`define MP2_3_PINCTRL_0_OD 0
`define MP2_3_PULLEN 0
`define MP2_3_PULLSEL 0
`define MP2_3_pad_y 0
`define MP2_4 0
`define MP2_4_GPIO_OUTPUT_ENABLE 0
`define MP2_4_INFUNC_EN 0
`define MP2_4_OUTFUNC_SEL 0
`define MP2_4_PINCTRL_0_IE 0
`define MP2_4_PINCTRL_0_OD 0
`define MP2_4_PULLEN 0
`define MP2_4_PULLSEL 0
`define MP2_4_pad_y 0
`define MP2_5 0
`define MP2_5_GPIO_OUTPUT_ENABLE 0
`define MP2_5_INFUNC_EN 0
`define MP2_5_OUTFUNC_SEL 0
`define MP2_5_PINCTRL_0_IE 0
`define MP2_5_PINCTRL_0_OD 0
`define MP2_5_PULLEN 0
`define MP2_5_PULLSEL 0
`define MP2_5_pad_y 0
`define MP2_6 0
`define MP2_6_GPIO_OUTPUT_ENABLE 0
`define MP2_6_INFUNC_EN 0
`define MP2_6_OUTFUNC_SEL 0
`define MP2_6_PINCTRL_0_IE 0
`define MP2_6_PINCTRL_0_OD 0
`define MP2_6_PULLEN 0
`define MP2_6_PULLSEL 0
`define MP2_6_pad_y 0
`define MP2_7 0
`define MP2_7_GPIO_OUTPUT_ENABLE 0
`define MP2_7_INFUNC_EN 0
`define MP2_7_OUTFUNC_SEL 0
`define MP2_7_PINCTRL_0_IE 0
`define MP2_7_PINCTRL_0_OD 0
`define MP2_7_PULLEN 0
`define MP2_7_PULLSEL 0
`define MP2_7_pad_y 0
`define MP2_8 0
`define MP2_8_GPIO_OUTPUT_ENABLE 0
`define MP2_8_INFUNC_EN 0
`define MP2_8_OUTFUNC_SEL 0
`define MP2_8_PINCTRL_0_IE 0
`define MP2_8_PINCTRL_0_OD 0
`define MP2_8_PULLEN 0
`define MP2_8_PULLSEL 0
`define MP2_8_pad_y 0
`define MP2_9 0
`define MP2_9_GPIO_OUTPUT_ENABLE 0
`define MP2_9_INFUNC_EN 0
`define MP2_9_OUTFUNC_SEL 0
`define MP2_9_PINCTRL_0_IE 0
`define MP2_9_PINCTRL_0_OD 0
`define MP2_9_PULLEN 0
`define MP2_9_PULLSEL 0
`define MP2_9_pad_y 0
`define MSC0CLK_IN 0
`define MSC0CLK_OE 0
`define MSC0CLK_OUT 0
`define MSC0CS0_IN 0
`define MSC0CS0_OE 0
`define MSC0CS0_OUT 0
`define MSC0CS1_IN 0
`define MSC0CS1_OE 0
`define MSC0CS1_OUT 0
`define MSC0CS2_IN 0
`define MSC0CS2_OE 0
`define MSC0CS2_OUT 0
`define MSC0CS3_IN 0
`define MSC0CS3_OE 0
`define MSC0CS3_OUT 0
`define MSC0SI_IN 0
`define MSC0SI_OE 0
`define MSC0SI_OUT 0
`define MSC0SO_IN 0
`define MSC0SO_OE 0
`define MSC0SO_OUT 0
`define MSC1CLK_IN 0
`define MSC1CLK_OE 0
`define MSC1CLK_OUT 0
`define MSC1CS0_IN 0
`define MSC1CS0_OE 0
`define MSC1CS0_OUT 0
`define MSC1CS1_IN 0
`define MSC1CS1_OE 0
`define MSC1CS1_OUT 0
`define MSC1CS2_IN 0
`define MSC1CS2_OE 0
`define MSC1CS2_OUT 0
`define MSC1CS3_IN 0
`define MSC1CS3_OE 0
`define MSC1CS3_OUT 0
`define MSC1SI_IN 0
`define MSC1SI_OE 0
`define MSC1SI_OUT 0
`define MSC1SO_IN 0
`define MSC1SO_OE 0
`define MSC1SO_OUT 0
`define OUTPUTXBAR0_IN 0
`define OUTPUTXBAR0_OE 0
`define OUTPUTXBAR0_OUT 0
`define OUTPUTXBAR10_IN 0
`define OUTPUTXBAR10_OE 0
`define OUTPUTXBAR10_OUT 0
`define OUTPUTXBAR11_IN 0
`define OUTPUTXBAR11_OE 0
`define OUTPUTXBAR11_OUT 0
`define OUTPUTXBAR12_IN 0
`define OUTPUTXBAR12_OE 0
`define OUTPUTXBAR12_OUT 0
`define OUTPUTXBAR13_IN 0
`define OUTPUTXBAR13_OE 0
`define OUTPUTXBAR13_OUT 0
`define OUTPUTXBAR14_IN 0
`define OUTPUTXBAR14_OE 0
`define OUTPUTXBAR14_OUT 0
`define OUTPUTXBAR15_IN 0
`define OUTPUTXBAR15_OE 0
`define OUTPUTXBAR15_OUT 0
`define OUTPUTXBAR1_IN 0
`define OUTPUTXBAR1_OE 0
`define OUTPUTXBAR1_OUT 0
`define OUTPUTXBAR2_IN 0
`define OUTPUTXBAR2_OE 0
`define OUTPUTXBAR2_OUT 0
`define OUTPUTXBAR3_IN 0
`define OUTPUTXBAR3_OE 0
`define OUTPUTXBAR3_OUT 0
`define OUTPUTXBAR4_IN 0
`define OUTPUTXBAR4_OE 0
`define OUTPUTXBAR4_OUT 0
`define OUTPUTXBAR5_IN 0
`define OUTPUTXBAR5_OE 0
`define OUTPUTXBAR5_OUT 0
`define OUTPUTXBAR6_IN 0
`define OUTPUTXBAR6_OE 0
`define OUTPUTXBAR6_OUT 0
`define OUTPUTXBAR7_IN 0
`define OUTPUTXBAR7_OE 0
`define OUTPUTXBAR7_OUT 0
`define OUTPUTXBAR8_IN 0
`define OUTPUTXBAR8_OE 0
`define OUTPUTXBAR8_OUT 0
`define OUTPUTXBAR9_IN 0
`define OUTPUTXBAR9_OE 0
`define OUTPUTXBAR9_OUT 0
`define PSI5_0_RX_IN 0
`define PSI5_0_RX_OE 0
`define PSI5_0_RX_OUT 0
`define PSI5_0_TX_IN 0
`define PSI5_0_TX_OE 0
`define PSI5_0_TX_OUT 0
`define PSI5_1_RX_IN 0
`define PSI5_1_RX_OE 0
`define PSI5_1_RX_OUT 0
`define PSI5_1_TX_IN 0
`define PSI5_1_TX_OE 0
`define PSI5_1_TX_OUT 0
`define PSI5_2_RX_IN 0
`define PSI5_2_RX_OE 0
`define PSI5_2_RX_OUT 0
`define PSI5_2_TX_IN 0
`define PSI5_2_TX_OE 0
`define PSI5_2_TX_OUT 0
`define PSI5_3_RX_IN 0
`define PSI5_3_RX_OE 0
`define PSI5_3_RX_OUT 0
`define PSI5_3_TX_IN 0
`define PSI5_3_TX_OE 0
`define PSI5_3_TX_OUT 0
`define PULL_DOWN 0
`define PULL_UP 1
`define RDC0PWM_N_IN 0
`define RDC0PWM_N_OE 0
`define RDC0PWM_N_OUT 0
`define RDC0PWM_P_IN 0
`define RDC0PWM_P_OE 0
`define RDC0PWM_P_OUT 0
`define RDC1PWM_N_IN 0
`define RDC1PWM_N_OE 0
`define RDC1PWM_N_OUT 0
`define RDC1PWM_P_IN 0
`define RDC1PWM_P_OE 0
`define RDC1PWM_P_OUT 0
`define RGMII0RXCLK_IN 0
`define RGMII0RXCLK_OE 0
`define RGMII0RXCLK_OUT 0
`define RGMII0RXCTL_IN 0
`define RGMII0RXCTL_OE 0
`define RGMII0RXCTL_OUT 0
`define RGMII0RXD0_IN 0
`define RGMII0RXD0_OE 0
`define RGMII0RXD0_OUT 0
`define RGMII0RXD1_IN 0
`define RGMII0RXD1_OE 0
`define RGMII0RXD1_OUT 0
`define RGMII0RXD2_IN 0
`define RGMII0RXD2_OE 0
`define RGMII0RXD2_OUT 0
`define RGMII0RXD3_IN 0
`define RGMII0RXD3_OE 0
`define RGMII0RXD3_OUT 0
`define RGMII0TXCLK_IN 0
`define RGMII0TXCLK_OE 0
`define RGMII0TXCLK_OUT 0
`define RGMII0TXCTL_IN 0
`define RGMII0TXCTL_OE 0
`define RGMII0TXCTL_OUT 0
`define RGMII0TXD0_IN 0
`define RGMII0TXD0_OE 0
`define RGMII0TXD0_OUT 0
`define RGMII0TXD1_IN 0
`define RGMII0TXD1_OE 0
`define RGMII0TXD1_OUT 0
`define RGMII0TXD2_IN 0
`define RGMII0TXD2_OE 0
`define RGMII0TXD2_OUT 0
`define RGMII0TXD3_IN 0
`define RGMII0TXD3_OE 0
`define RGMII0TXD3_OUT 0
`define RGMII1RXCLK_IN 0
`define RGMII1RXCLK_OE 0
`define RGMII1RXCLK_OUT 0
`define RGMII1RXCTL_IN 0
`define RGMII1RXCTL_OE 0
`define RGMII1RXCTL_OUT 0
`define RGMII1RXD0_IN 0
`define RGMII1RXD0_OE 0
`define RGMII1RXD0_OUT 0
`define RGMII1RXD1_IN 0
`define RGMII1RXD1_OE 0
`define RGMII1RXD1_OUT 0
`define RGMII1RXD2_IN 0
`define RGMII1RXD2_OE 0
`define RGMII1RXD2_OUT 0
`define RGMII1RXD3_IN 0
`define RGMII1RXD3_OE 0
`define RGMII1RXD3_OUT 0
`define RGMII1TXCLK_IN 0
`define RGMII1TXCLK_OE 0
`define RGMII1TXCLK_OUT 0
`define RGMII1TXCTL_IN 0
`define RGMII1TXCTL_OE 0
`define RGMII1TXCTL_OUT 0
`define RGMII1TXD0_IN 0
`define RGMII1TXD0_OE 0
`define RGMII1TXD0_OUT 0
`define RGMII1TXD1_IN 0
`define RGMII1TXD1_OE 0
`define RGMII1TXD1_OUT 0
`define RGMII1TXD2_IN 0
`define RGMII1TXD2_OE 0
`define RGMII1TXD2_OUT 0
`define RGMII1TXD3_IN 0
`define RGMII1TXD3_OE 0
`define RGMII1TXD3_OUT 0
`define RGMII2RXCLK_IN 0
`define RGMII2RXCLK_OE 0
`define RGMII2RXCLK_OUT 0
`define RGMII2RXCTL_IN 0
`define RGMII2RXCTL_OE 0
`define RGMII2RXCTL_OUT 0
`define RGMII2RXD0_IN 0
`define RGMII2RXD0_OE 0
`define RGMII2RXD0_OUT 0
`define RGMII2RXD1_IN 0
`define RGMII2RXD1_OE 0
`define RGMII2RXD1_OUT 0
`define RGMII2RXD2_IN 0
`define RGMII2RXD2_OE 0
`define RGMII2RXD2_OUT 0
`define RGMII2RXD3_IN 0
`define RGMII2RXD3_OE 0
`define RGMII2RXD3_OUT 0
`define RGMII2TXCLK_IN 0
`define RGMII2TXCLK_OE 0
`define RGMII2TXCLK_OUT 0
`define RGMII2TXCTL_IN 0
`define RGMII2TXCTL_OE 0
`define RGMII2TXCTL_OUT 0
`define RGMII2TXD0_IN 0
`define RGMII2TXD0_OE 0
`define RGMII2TXD0_OUT 0
`define RGMII2TXD1_IN 0
`define RGMII2TXD1_OE 0
`define RGMII2TXD1_OUT 0
`define RGMII2TXD2_IN 0
`define RGMII2TXD2_OE 0
`define RGMII2TXD2_OUT 0
`define RGMII2TXD3_IN 0
`define RGMII2TXD3_OE 0
`define RGMII2TXD3_OUT 0
`define SDFM0CLK_IN 0
`define SDFM0DATA_IN 0
`define SDFM10CLK_IN 0
`define SDFM10DATA_IN 0
`define SDFM11CLK_IN 0
`define SDFM11DATA_IN 0
`define SDFM1CLK_IN 0
`define SDFM1DATA_IN 0
`define SDFM2CLK_IN 0
`define SDFM2DATA_IN 0
`define SDFM3CLK_IN 0
`define SDFM3DATA_IN 0
`define SDFM4CLK_IN 0
`define SDFM4DATA_IN 0
`define SDFM5CLK_IN 0
`define SDFM5DATA_IN 0
`define SDFM6CLK_IN 0
`define SDFM6DATA_IN 0
`define SDFM7CLK_IN 0
`define SDFM7DATA_IN 0
`define SDFM8CLK_IN 0
`define SDFM8DATA_IN 0
`define SDFM9CLK_IN 0
`define SDFM9DATA_IN 0
`define SENT0TXRX_IN 0
`define SENT0TXRX_OE 0
`define SENT0TXRX_OUT 0
`define SENT1TXRX_IN 0
`define SENT1TXRX_OE 0
`define SENT1TXRX_OUT 0
`define SENT2TXRX_IN 0
`define SENT2TXRX_OE 0
`define SENT2TXRX_OUT 0
`define SENT3TXRX_IN 0
`define SENT3TXRX_OE 0
`define SENT3TXRX_OUT 0
`define SENT4TXRX_IN 0
`define SENT4TXRX_OE 0
`define SENT4TXRX_OUT 0
`define SENT5TXRX_IN 0
`define SENT5TXRX_OE 0
`define SENT5TXRX_OUT 0
`define SPI2CLK_IN 0
`define SPI2CLK_OE 0
`define SPI2CLK_OUT 0
`define SPI2CS0_IN 0
`define SPI2CS0_OE 0
`define SPI2CS0_OUT 0
`define SPI2CS1_IN 0
`define SPI2CS1_OE 0
`define SPI2CS1_OUT 0
`define SPI2CS2_IN 0
`define SPI2CS2_OE 0
`define SPI2CS2_OUT 0
`define SPI2CS3_IN 0
`define SPI2CS3_OE 0
`define SPI2CS3_OUT 0
`define SPI2CS4_IN 0
`define SPI2CS4_OE 0
`define SPI2CS4_OUT 0
`define SPI2CS5_IN 0
`define SPI2CS5_OE 0
`define SPI2CS5_OUT 0
`define SPI2PICO_IN 0
`define SPI2PICO_OE 0
`define SPI2PICO_OUT 0
`define SPI2POCI_IN 0
`define SPI2POCI_OE 0
`define SPI2POCI_OUT 0
`define SPI3CLK_IN 0
`define SPI3CLK_OE 0
`define SPI3CLK_OUT 0
`define SPI3CS0_IN 0
`define SPI3CS0_OE 0
`define SPI3CS0_OUT 0
`define SPI3CS1_IN 0
`define SPI3CS1_OE 0
`define SPI3CS1_OUT 0
`define SPI3CS2_IN 0
`define SPI3CS2_OE 0
`define SPI3CS2_OUT 0
`define SPI3CS3_IN 0
`define SPI3CS3_OE 0
`define SPI3CS3_OUT 0
`define SPI3CS4_IN 0
`define SPI3CS4_OE 0
`define SPI3CS4_OUT 0
`define SPI3CS5_IN 0
`define SPI3CS5_OE 0
`define SPI3CS5_OUT 0
`define SPI3PICO_IN 0
`define SPI3PICO_OE 0
`define SPI3PICO_OUT 0
`define SPI3POCI_IN 0
`define SPI3POCI_OE 0
`define SPI3POCI_OUT 0
`define SPI4CLK_IN 0
`define SPI4CLK_OE 0
`define SPI4CLK_OUT 0
`define SPI4CS0_IN 0
`define SPI4CS0_OE 0
`define SPI4CS0_OUT 0
`define SPI4CS1_IN 0
`define SPI4CS1_OE 0
`define SPI4CS1_OUT 0
`define SPI4CS2_IN 0
`define SPI4CS2_OE 0
`define SPI4CS2_OUT 0
`define SPI4CS3_IN 0
`define SPI4CS3_OE 0
`define SPI4CS3_OUT 0
`define SPI4CS4_IN 0
`define SPI4CS4_OE 0
`define SPI4CS4_OUT 0
`define SPI4CS5_IN 0
`define SPI4CS5_OE 0
`define SPI4CS5_OUT 0
`define SPI4PICO_IN 0
`define SPI4PICO_OE 0
`define SPI4PICO_OUT 0
`define SPI4POCI_IN 0
`define SPI4POCI_OE 0
`define SPI4POCI_OUT 0
`define SPI5CLK_IN 0
`define SPI5CLK_OE 0
`define SPI5CLK_OUT 0
`define SPI5CS0_IN 0
`define SPI5CS0_OE 0
`define SPI5CS0_OUT 0
`define SPI5CS1_IN 0
`define SPI5CS1_OE 0
`define SPI5CS1_OUT 0
`define SPI5CS2_IN 0
`define SPI5CS2_OE 0
`define SPI5CS2_OUT 0
`define SPI5CS3_IN 0
`define SPI5CS3_OE 0
`define SPI5CS3_OUT 0
`define SPI5CS4_IN 0
`define SPI5CS4_OE 0
`define SPI5CS4_OUT 0
`define SPI5CS5_IN 0
`define SPI5CS5_OE 0
`define SPI5CS5_OUT 0
`define SPI5PICO_IN 0
`define SPI5PICO_OE 0
`define SPI5PICO_OUT 0
`define SPI5POCI_IN 0
`define SPI5POCI_OE 0
`define SPI5POCI_OUT 0
`define SPI6CLK_IN 0
`define SPI6CLK_OE 0
`define SPI6CLK_OUT 0
`define SPI6CS0_IN 0
`define SPI6CS0_OE 0
`define SPI6CS0_OUT 0
`define SPI6CS1_IN 0
`define SPI6CS1_OE 0
`define SPI6CS1_OUT 0
`define SPI6CS2_IN 0
`define SPI6CS2_OE 0
`define SPI6CS2_OUT 0
`define SPI6CS3_IN 0
`define SPI6CS3_OE 0
`define SPI6CS3_OUT 0
`define SPI6CS4_IN 0
`define SPI6CS4_OE 0
`define SPI6CS4_OUT 0
`define SPI6CS5_IN 0
`define SPI6CS5_OE 0
`define SPI6CS5_OUT 0
`define SPI6PICO_IN 0
`define SPI6PICO_OE 0
`define SPI6PICO_OUT 0
`define SPI6POCI_IN 0
`define SPI6POCI_OE 0
`define SPI6POCI_OUT 0
`define SPI7CLK_IN 0
`define SPI7CLK_OE 0
`define SPI7CLK_OUT 0
`define SPI7CS0_IN 0
`define SPI7CS0_OE 0
`define SPI7CS0_OUT 0
`define SPI7CS1_IN 0
`define SPI7CS1_OE 0
`define SPI7CS1_OUT 0
`define SPI7CS2_IN 0
`define SPI7CS2_OE 0
`define SPI7CS2_OUT 0
`define SPI7CS3_IN 0
`define SPI7CS3_OE 0
`define SPI7CS3_OUT 0
`define SPI7CS4_IN 0
`define SPI7CS4_OE 0
`define SPI7CS4_OUT 0
`define SPI7CS5_IN 0
`define SPI7CS5_OE 0
`define SPI7CS5_OUT 0
`define SPI7PICO_IN 0
`define SPI7PICO_OE 0
`define SPI7PICO_OUT 0
`define SPI7POCI_IN 0
`define SPI7POCI_OE 0
`define SPI7POCI_OUT 0
`define SPI8CLK_IN 0
`define SPI8CLK_OE 0
`define SPI8CLK_OUT 0
`define SPI8CS0_IN 0
`define SPI8CS0_OE 0
`define SPI8CS0_OUT 0
`define SPI8CS1_IN 0
`define SPI8CS1_OE 0
`define SPI8CS1_OUT 0
`define SPI8CS2_IN 0
`define SPI8CS2_OE 0
`define SPI8CS2_OUT 0
`define SPI8CS3_IN 0
`define SPI8CS3_OE 0
`define SPI8CS3_OUT 0
`define SPI8CS4_IN 0
`define SPI8CS4_OE 0
`define SPI8CS4_OUT 0
`define SPI8CS5_IN 0
`define SPI8CS5_OE 0
`define SPI8CS5_OUT 0
`define SPI8PICO_IN 0
`define SPI8PICO_OE 0
`define SPI8PICO_OUT 0
`define SPI8POCI_IN 0
`define SPI8POCI_OE 0
`define SPI8POCI_OUT 0
`define SPI9CLK_IN 0
`define SPI9CLK_OE 0
`define SPI9CLK_OUT 0
`define SPI9CS0_IN 0
`define SPI9CS0_OE 0
`define SPI9CS0_OUT 0
`define SPI9CS1_IN 0
`define SPI9CS1_OE 0
`define SPI9CS1_OUT 0
`define SPI9CS2_IN 0
`define SPI9CS2_OE 0
`define SPI9CS2_OUT 0
`define SPI9CS3_IN 0
`define SPI9CS3_OE 0
`define SPI9CS3_OUT 0
`define SPI9CS4_IN 0
`define SPI9CS4_OE 0
`define SPI9CS4_OUT 0
`define SPI9CS5_IN 0
`define SPI9CS5_OE 0
`define SPI9CS5_OUT 0
`define SPI9PICO_IN 0
`define SPI9PICO_OE 0
`define SPI9PICO_OUT 0
`define SPI9POCI_IN 0
`define SPI9POCI_OE 0
`define SPI9POCI_OUT 0
`define T1S0ED_IN 0
`define T1S0ED_OE 0
`define T1S0ED_OUT 0
`define T1S0RX_IN 0
`define T1S0RX_OE 0
`define T1S0RX_OUT 0
`define T1S0TX_IN 0
`define T1S0TX_OE 0
`define T1S0TX_OUT 0
`define T1S1ED_IN 0
`define T1S1ED_OE 0
`define T1S1ED_OUT 0
`define T1S1RX_IN 0
`define T1S1RX_OE 0
`define T1S1RX_OUT 0
`define T1S1TX_IN 0
`define T1S1TX_OE 0
`define T1S1TX_OUT 0
`define T1S2ED_IN 0
`define T1S2ED_OE 0
`define T1S2ED_OUT 0
`define T1S2RX_IN 0
`define T1S2RX_OE 0
`define T1S2RX_OUT 0
`define T1S2TX_IN 0
`define T1S2TX_OE 0
`define T1S2TX_OUT 0
`define T1S3ED_IN 0
`define T1S3ED_OE 0
`define T1S3ED_OUT 0
`define T1S3RX_IN 0
`define T1S3RX_OE 0
`define T1S3RX_OUT 0
`define T1S3TX_IN 0
`define T1S3TX_OE 0
`define T1S3TX_OUT 0
`define T1SMDC_IN 0
`define T1SMDC_OE 0
`define T1SMDC_OUT 0
`define T1SMDIO_IN 0
`define T1SMDIO_OE 0
`define T1SMDIO_OUT 0
`define TPIUCLK_IN 0
`define TPIUCLK_OE 0
`define TPIUCLK_OUT 0
`define TPIUCTL_IN 0
`define TPIUCTL_OE 0
`define TPIUCTL_OUT 0
`define TPIUDATA0_IN 0
`define TPIUDATA0_OE 0
`define TPIUDATA0_OUT 0
`define TPIUDATA1_IN 0
`define TPIUDATA1_OE 0
`define TPIUDATA1_OUT 0
`define TPIUDATA2_IN 0
`define TPIUDATA2_OE 0
`define TPIUDATA2_OUT 0
`define TPIUDATA3_IN 0
`define TPIUDATA3_OE 0
`define TPIUDATA3_OUT 0
`define UART0RX_IN 0
`define UART0RX_OE 0
`define UART0RX_OUT 0
`define UART0TX_IN 0
`define UART0TX_OE 0
`define UART0TX_OUT 0
`define UART1RX_IN 0
`define UART1RX_OE 0
`define UART1RX_OUT 0
`define UART1TX_IN 0
`define UART1TX_OE 0
`define UART1TX_OUT 0
`define XSPI0CLK_IN 0
`define XSPI0CLK_OE 0
`define XSPI0CLK_OUT 0
`define XSPI0CS0_IN 0
`define XSPI0CS0_OE 0
`define XSPI0CS0_OUT 0
`define XSPI0CS1_IN 0
`define XSPI0CS1_OE 0
`define XSPI0CS1_OUT 0
`define XSPI0DQS_IN 0
`define XSPI0DQS_OE 0
`define XSPI0DQS_OUT 0
`define XSPI0DS0_IN 0
`define XSPI0DS0_OE 0
`define XSPI0DS0_OUT 0
`define XSPI0DS1_IN 0
`define XSPI0DS1_OE 0
`define XSPI0DS1_OUT 0
`define XSPI0DS2_IN 0
`define XSPI0DS2_OE 0
`define XSPI0DS2_OUT 0
`define XSPI0DS3_IN 0
`define XSPI0DS3_OE 0
`define XSPI0DS3_OUT 0
`define XSPI0DS4_IN 0
`define XSPI0DS4_OE 0
`define XSPI0DS4_OUT 0
`define XSPI0DS5_IN 0
`define XSPI0DS5_OE 0
`define XSPI0DS5_OUT 0
`define XSPI0DS6_IN 0
`define XSPI0DS6_OE 0
`define XSPI0DS6_OUT 0
`define XSPI0DS7_IN 0
`define XSPI0DS7_OE 0
`define XSPI0DS7_OUT 0
`define default_value 0
`define input_func_concat_DP0_0 0
`define input_func_concat_DP0_1 0
`define input_func_concat_DP0_10 0
`define input_func_concat_DP0_11 0
`define input_func_concat_DP0_12 0
`define input_func_concat_DP0_13 0
`define input_func_concat_DP0_14 0
`define input_func_concat_DP0_15 0
`define input_func_concat_DP0_16 0
`define input_func_concat_DP0_17 0
`define input_func_concat_DP0_18 0
`define input_func_concat_DP0_19 0
`define input_func_concat_DP0_2 0
`define input_func_concat_DP0_20 0
`define input_func_concat_DP0_21 0
`define input_func_concat_DP0_22 0
`define input_func_concat_DP0_23 0
`define input_func_concat_DP0_24 0
`define input_func_concat_DP0_25 0
`define input_func_concat_DP0_26 0
`define input_func_concat_DP0_27 0
`define input_func_concat_DP0_28 0
`define input_func_concat_DP0_29 0
`define input_func_concat_DP0_3 0
`define input_func_concat_DP0_30 0
`define input_func_concat_DP0_31 0
`define input_func_concat_DP0_4 0
`define input_func_concat_DP0_5 0
`define input_func_concat_DP0_6 0
`define input_func_concat_DP0_7 0
`define input_func_concat_DP0_8 0
`define input_func_concat_DP0_9 0
`define input_func_concat_DP1_0 0
`define input_func_concat_DP1_1 0
`define input_func_concat_DP1_10 0
`define input_func_concat_DP1_11 0
`define input_func_concat_DP1_12 0
`define input_func_concat_DP1_13 0
`define input_func_concat_DP1_14 0
`define input_func_concat_DP1_15 0
`define input_func_concat_DP1_16 0
`define input_func_concat_DP1_17 0
`define input_func_concat_DP1_18 0
`define input_func_concat_DP1_19 0
`define input_func_concat_DP1_2 0
`define input_func_concat_DP1_20 0
`define input_func_concat_DP1_21 0
`define input_func_concat_DP1_22 0
`define input_func_concat_DP1_23 0
`define input_func_concat_DP1_24 0
`define input_func_concat_DP1_25 0
`define input_func_concat_DP1_26 0
`define input_func_concat_DP1_27 0
`define input_func_concat_DP1_28 0
`define input_func_concat_DP1_29 0
`define input_func_concat_DP1_3 0
`define input_func_concat_DP1_30 0
`define input_func_concat_DP1_31 0
`define input_func_concat_DP1_4 0
`define input_func_concat_DP1_5 0
`define input_func_concat_DP1_6 0
`define input_func_concat_DP1_7 0
`define input_func_concat_DP1_8 0
`define input_func_concat_DP1_9 0
`define input_func_concat_DP2_0 0
`define input_func_concat_DP2_1 0
`define input_func_concat_DP2_10 0
`define input_func_concat_DP2_11 0
`define input_func_concat_DP2_12 0
`define input_func_concat_DP2_13 0
`define input_func_concat_DP2_14 0
`define input_func_concat_DP2_15 0
`define input_func_concat_DP2_16 0
`define input_func_concat_DP2_17 0
`define input_func_concat_DP2_18 0
`define input_func_concat_DP2_19 0
`define input_func_concat_DP2_2 0
`define input_func_concat_DP2_20 0
`define input_func_concat_DP2_21 0
`define input_func_concat_DP2_22 0
`define input_func_concat_DP2_23 0
`define input_func_concat_DP2_24 0
`define input_func_concat_DP2_25 0
`define input_func_concat_DP2_26 0
`define input_func_concat_DP2_27 0
`define input_func_concat_DP2_28 0
`define input_func_concat_DP2_29 0
`define input_func_concat_DP2_3 0
`define input_func_concat_DP2_30 0
`define input_func_concat_DP2_31 0
`define input_func_concat_DP2_4 0
`define input_func_concat_DP2_5 0
`define input_func_concat_DP2_6 0
`define input_func_concat_DP2_7 0
`define input_func_concat_DP2_8 0
`define input_func_concat_DP2_9 0
`define input_func_concat_DP3_0 0
`define input_func_concat_DP3_1 0
`define input_func_concat_DP3_10 0
`define input_func_concat_DP3_11 0
`define input_func_concat_DP3_12 0
`define input_func_concat_DP3_13 0
`define input_func_concat_DP3_14 0
`define input_func_concat_DP3_15 0
`define input_func_concat_DP3_16 0
`define input_func_concat_DP3_17 0
`define input_func_concat_DP3_18 0
`define input_func_concat_DP3_19 0
`define input_func_concat_DP3_2 0
`define input_func_concat_DP3_20 0
`define input_func_concat_DP3_21 0
`define input_func_concat_DP3_22 0
`define input_func_concat_DP3_23 0
`define input_func_concat_DP3_24 0
`define input_func_concat_DP3_25 0
`define input_func_concat_DP3_26 0
`define input_func_concat_DP3_27 0
`define input_func_concat_DP3_28 0
`define input_func_concat_DP3_29 0
`define input_func_concat_DP3_3 0
`define input_func_concat_DP3_30 0
`define input_func_concat_DP3_31 0
`define input_func_concat_DP3_4 0
`define input_func_concat_DP3_5 0
`define input_func_concat_DP3_6 0
`define input_func_concat_DP3_7 0
`define input_func_concat_DP3_8 0
`define input_func_concat_DP3_9 0
`define input_func_concat_DP4_0 0
`define input_func_concat_DP4_1 0
`define input_func_concat_DP4_10 0
`define input_func_concat_DP4_11 0
`define input_func_concat_DP4_12 0
`define input_func_concat_DP4_13 0
`define input_func_concat_DP4_14 0
`define input_func_concat_DP4_15 0
`define input_func_concat_DP4_16 0
`define input_func_concat_DP4_17 0
`define input_func_concat_DP4_18 0
`define input_func_concat_DP4_19 0
`define input_func_concat_DP4_2 0
`define input_func_concat_DP4_20 0
`define input_func_concat_DP4_21 0
`define input_func_concat_DP4_22 0
`define input_func_concat_DP4_23 0
`define input_func_concat_DP4_24 0
`define input_func_concat_DP4_25 0
`define input_func_concat_DP4_26 0
`define input_func_concat_DP4_27 0
`define input_func_concat_DP4_28 0
`define input_func_concat_DP4_29 0
`define input_func_concat_DP4_3 0
`define input_func_concat_DP4_30 0
`define input_func_concat_DP4_31 0
`define input_func_concat_DP4_4 0
`define input_func_concat_DP4_5 0
`define input_func_concat_DP4_6 0
`define input_func_concat_DP4_7 0
`define input_func_concat_DP4_8 0
`define input_func_concat_DP4_9 0
`define input_func_concat_DP5_0 0
`define input_func_concat_DP5_1 0
`define input_func_concat_DP5_10 0
`define input_func_concat_DP5_11 0
`define input_func_concat_DP5_12 0
`define input_func_concat_DP5_13 0
`define input_func_concat_DP5_14 0
`define input_func_concat_DP5_15 0
`define input_func_concat_DP5_16 0
`define input_func_concat_DP5_17 0
`define input_func_concat_DP5_18 0
`define input_func_concat_DP5_19 0
`define input_func_concat_DP5_2 0
`define input_func_concat_DP5_20 0
`define input_func_concat_DP5_21 0
`define input_func_concat_DP5_22 0
`define input_func_concat_DP5_23 0
`define input_func_concat_DP5_24 0
`define input_func_concat_DP5_25 0
`define input_func_concat_DP5_26 0
`define input_func_concat_DP5_27 0
`define input_func_concat_DP5_28 0
`define input_func_concat_DP5_29 0
`define input_func_concat_DP5_3 0
`define input_func_concat_DP5_30 0
`define input_func_concat_DP5_31 0
`define input_func_concat_DP5_4 0
`define input_func_concat_DP5_5 0
`define input_func_concat_DP5_6 0
`define input_func_concat_DP5_7 0
`define input_func_concat_DP5_8 0
`define input_func_concat_DP5_9 0
`define input_func_concat_DP6_0 0
`define input_func_concat_DP6_1 0
`define input_func_concat_DP6_10 0
`define input_func_concat_DP6_11 0
`define input_func_concat_DP6_12 0
`define input_func_concat_DP6_13 0
`define input_func_concat_DP6_14 0
`define input_func_concat_DP6_15 0
`define input_func_concat_DP6_16 0
`define input_func_concat_DP6_17 0
`define input_func_concat_DP6_18 0
`define input_func_concat_DP6_19 0
`define input_func_concat_DP6_2 0
`define input_func_concat_DP6_20 0
`define input_func_concat_DP6_21 0
`define input_func_concat_DP6_22 0
`define input_func_concat_DP6_23 0
`define input_func_concat_DP6_24 0
`define input_func_concat_DP6_25 0
`define input_func_concat_DP6_26 0
`define input_func_concat_DP6_27 0
`define input_func_concat_DP6_3 0
`define input_func_concat_DP6_4 0
`define input_func_concat_DP6_5 0
`define input_func_concat_DP6_6 0
`define input_func_concat_DP6_7 0
`define input_func_concat_DP6_8 0
`define input_func_concat_DP6_9 0
`define input_func_concat_DP7_0 0
`define input_func_concat_DP7_1 0
`define input_func_concat_DP7_10 0
`define input_func_concat_DP7_11 0
`define input_func_concat_DP7_12 0
`define input_func_concat_DP7_13 0
`define input_func_concat_DP7_14 0
`define input_func_concat_DP7_15 0
`define input_func_concat_DP7_2 0
`define input_func_concat_DP7_3 0
`define input_func_concat_DP7_4 0
`define input_func_concat_DP7_5 0
`define input_func_concat_DP7_6 0
`define input_func_concat_DP7_7 0
`define input_func_concat_DP7_8 0
`define input_func_concat_DP7_9 0
`define input_func_concat_MP0_0 0
`define input_func_concat_MP0_1 0
`define input_func_concat_MP0_10 0
`define input_func_concat_MP0_11 0
`define input_func_concat_MP0_12 0
`define input_func_concat_MP0_13 0
`define input_func_concat_MP0_14 0
`define input_func_concat_MP0_15 0
`define input_func_concat_MP0_16 0
`define input_func_concat_MP0_17 0
`define input_func_concat_MP0_18 0
`define input_func_concat_MP0_19 0
`define input_func_concat_MP0_2 0
`define input_func_concat_MP0_20 0
`define input_func_concat_MP0_21 0
`define input_func_concat_MP0_22 0
`define input_func_concat_MP0_23 0
`define input_func_concat_MP0_24 0
`define input_func_concat_MP0_25 0
`define input_func_concat_MP0_26 0
`define input_func_concat_MP0_27 0
`define input_func_concat_MP0_28 0
`define input_func_concat_MP0_29 0
`define input_func_concat_MP0_3 0
`define input_func_concat_MP0_30 0
`define input_func_concat_MP0_31 0
`define input_func_concat_MP0_4 0
`define input_func_concat_MP0_5 0
`define input_func_concat_MP0_6 0
`define input_func_concat_MP0_7 0
`define input_func_concat_MP0_8 0
`define input_func_concat_MP0_9 0
`define input_func_concat_MP1_0 0
`define input_func_concat_MP1_1 0
`define input_func_concat_MP1_10 0
`define input_func_concat_MP1_11 0
`define input_func_concat_MP1_12 0
`define input_func_concat_MP1_13 0
`define input_func_concat_MP1_14 0
`define input_func_concat_MP1_15 0
`define input_func_concat_MP1_2 0
`define input_func_concat_MP1_3 0
`define input_func_concat_MP1_4 0
`define input_func_concat_MP1_5 0
`define input_func_concat_MP1_6 0
`define input_func_concat_MP1_7 0
`define input_func_concat_MP1_8 0
`define input_func_concat_MP1_9 0
`define input_func_concat_MP2_0 0
`define input_func_concat_MP2_1 0
`define input_func_concat_MP2_10 0
`define input_func_concat_MP2_11 0
`define input_func_concat_MP2_12 0
`define input_func_concat_MP2_13 0
`define input_func_concat_MP2_14 0
`define input_func_concat_MP2_15 0
`define input_func_concat_MP2_2 0
`define input_func_concat_MP2_3 0
`define input_func_concat_MP2_4 0
`define input_func_concat_MP2_5 0
`define input_func_concat_MP2_6 0
`define input_func_concat_MP2_7 0
`define input_func_concat_MP2_8 0
`define input_func_concat_MP2_9 0
`define nan_IN 0
wire [31:0] input_func_concat_DP0_0;
wire [31:0] input_func_concat_DP0_10;
wire [31:0] input_func_concat_DP0_11;
wire [31:0] input_func_concat_DP0_12;
wire [31:0] input_func_concat_DP0_13;
wire [31:0] input_func_concat_DP0_14;
wire [31:0] input_func_concat_DP0_15;
wire [31:0] input_func_concat_DP0_16;
wire [31:0] input_func_concat_DP0_17;
wire [31:0] input_func_concat_DP0_18;
wire [31:0] input_func_concat_DP0_19;
wire [31:0] input_func_concat_DP0_1;
wire [31:0] input_func_concat_DP0_20;
wire [31:0] input_func_concat_DP0_21;
wire [31:0] input_func_concat_DP0_22;
wire [31:0] input_func_concat_DP0_23;
wire [31:0] input_func_concat_DP0_24;
wire [31:0] input_func_concat_DP0_25;
wire [31:0] input_func_concat_DP0_26;
wire [31:0] input_func_concat_DP0_27;
wire [31:0] input_func_concat_DP0_28;
wire [31:0] input_func_concat_DP0_29;
wire [31:0] input_func_concat_DP0_2;
wire [31:0] input_func_concat_DP0_30;
wire [31:0] input_func_concat_DP0_31;
wire [31:0] input_func_concat_DP0_3;
wire [31:0] input_func_concat_DP0_4;
wire [31:0] input_func_concat_DP0_5;
wire [31:0] input_func_concat_DP0_6;
wire [31:0] input_func_concat_DP0_7;
wire [31:0] input_func_concat_DP0_8;
wire [31:0] input_func_concat_DP0_9;
wire [31:0] input_func_concat_DP1_0;
wire [31:0] input_func_concat_DP1_10;
wire [31:0] input_func_concat_DP1_11;
wire [31:0] input_func_concat_DP1_12;
wire [31:0] input_func_concat_DP1_13;
wire [31:0] input_func_concat_DP1_14;
wire [31:0] input_func_concat_DP1_15;
wire [31:0] input_func_concat_DP1_16;
wire [31:0] input_func_concat_DP1_17;
wire [31:0] input_func_concat_DP1_18;
wire [31:0] input_func_concat_DP1_19;
wire [31:0] input_func_concat_DP1_1;
wire [31:0] input_func_concat_DP1_20;
wire [31:0] input_func_concat_DP1_21;
wire [31:0] input_func_concat_DP1_22;
wire [31:0] input_func_concat_DP1_23;
wire [31:0] input_func_concat_DP1_24;
wire [31:0] input_func_concat_DP1_25;
wire [31:0] input_func_concat_DP1_26;
wire [31:0] input_func_concat_DP1_27;
wire [31:0] input_func_concat_DP1_28;
wire [31:0] input_func_concat_DP1_29;
wire [31:0] input_func_concat_DP1_2;
wire [31:0] input_func_concat_DP1_30;
wire [31:0] input_func_concat_DP1_31;
wire [31:0] input_func_concat_DP1_3;
wire [31:0] input_func_concat_DP1_4;
wire [31:0] input_func_concat_DP1_5;
wire [31:0] input_func_concat_DP1_6;
wire [31:0] input_func_concat_DP1_7;
wire [31:0] input_func_concat_DP1_8;
wire [31:0] input_func_concat_DP1_9;
wire [31:0] input_func_concat_DP2_0;
wire [31:0] input_func_concat_DP2_10;
wire [31:0] input_func_concat_DP2_11;
wire [31:0] input_func_concat_DP2_12;
wire [31:0] input_func_concat_DP2_13;
wire [31:0] input_func_concat_DP2_14;
wire [31:0] input_func_concat_DP2_15;
wire [31:0] input_func_concat_DP2_16;
wire [31:0] input_func_concat_DP2_17;
wire [31:0] input_func_concat_DP2_18;
wire [31:0] input_func_concat_DP2_19;
wire [31:0] input_func_concat_DP2_1;
wire [31:0] input_func_concat_DP2_20;
wire [31:0] input_func_concat_DP2_21;
wire [31:0] input_func_concat_DP2_22;
wire [31:0] input_func_concat_DP2_23;
wire [31:0] input_func_concat_DP2_24;
wire [31:0] input_func_concat_DP2_25;
wire [31:0] input_func_concat_DP2_26;
wire [31:0] input_func_concat_DP2_27;
wire [31:0] input_func_concat_DP2_28;
wire [31:0] input_func_concat_DP2_29;
wire [31:0] input_func_concat_DP2_2;
wire [31:0] input_func_concat_DP2_30;
wire [31:0] input_func_concat_DP2_31;
wire [31:0] input_func_concat_DP2_3;
wire [31:0] input_func_concat_DP2_4;
wire [31:0] input_func_concat_DP2_5;
wire [31:0] input_func_concat_DP2_6;
wire [31:0] input_func_concat_DP2_7;
wire [31:0] input_func_concat_DP2_8;
wire [31:0] input_func_concat_DP2_9;
wire [31:0] input_func_concat_DP3_0;
wire [31:0] input_func_concat_DP3_10;
wire [31:0] input_func_concat_DP3_11;
wire [31:0] input_func_concat_DP3_12;
wire [31:0] input_func_concat_DP3_13;
wire [31:0] input_func_concat_DP3_14;
wire [31:0] input_func_concat_DP3_15;
wire [31:0] input_func_concat_DP3_16;
wire [31:0] input_func_concat_DP3_17;
wire [31:0] input_func_concat_DP3_18;
wire [31:0] input_func_concat_DP3_19;
wire [31:0] input_func_concat_DP3_1;
wire [31:0] input_func_concat_DP3_20;
wire [31:0] input_func_concat_DP3_21;
wire [31:0] input_func_concat_DP3_22;
wire [31:0] input_func_concat_DP3_23;
wire [31:0] input_func_concat_DP3_24;
wire [31:0] input_func_concat_DP3_25;
wire [31:0] input_func_concat_DP3_26;
wire [31:0] input_func_concat_DP3_27;
wire [31:0] input_func_concat_DP3_28;
wire [31:0] input_func_concat_DP3_29;
wire [31:0] input_func_concat_DP3_2;
wire [31:0] input_func_concat_DP3_30;
wire [31:0] input_func_concat_DP3_31;
wire [31:0] input_func_concat_DP3_3;
wire [31:0] input_func_concat_DP3_4;
wire [31:0] input_func_concat_DP3_5;
wire [31:0] input_func_concat_DP3_6;
wire [31:0] input_func_concat_DP3_7;
wire [31:0] input_func_concat_DP3_8;
wire [31:0] input_func_concat_DP3_9;
wire [31:0] input_func_concat_DP4_0;
wire [31:0] input_func_concat_DP4_10;
wire [31:0] input_func_concat_DP4_11;
wire [31:0] input_func_concat_DP4_12;
wire [31:0] input_func_concat_DP4_13;
wire [31:0] input_func_concat_DP4_14;
wire [31:0] input_func_concat_DP4_15;
wire [31:0] input_func_concat_DP4_16;
wire [31:0] input_func_concat_DP4_17;
wire [31:0] input_func_concat_DP4_18;
wire [31:0] input_func_concat_DP4_19;
wire [31:0] input_func_concat_DP4_1;
wire [31:0] input_func_concat_DP4_20;
wire [31:0] input_func_concat_DP4_21;
wire [31:0] input_func_concat_DP4_22;
wire [31:0] input_func_concat_DP4_23;
wire [31:0] input_func_concat_DP4_24;
wire [31:0] input_func_concat_DP4_25;
wire [31:0] input_func_concat_DP4_26;
wire [31:0] input_func_concat_DP4_27;
wire [31:0] input_func_concat_DP4_28;
wire [31:0] input_func_concat_DP4_29;
wire [31:0] input_func_concat_DP4_2;
wire [31:0] input_func_concat_DP4_30;
wire [31:0] input_func_concat_DP4_31;
wire [31:0] input_func_concat_DP4_3;
wire [31:0] input_func_concat_DP4_4;
wire [31:0] input_func_concat_DP4_5;
wire [31:0] input_func_concat_DP4_6;
wire [31:0] input_func_concat_DP4_7;
wire [31:0] input_func_concat_DP4_8;
wire [31:0] input_func_concat_DP4_9;
wire [31:0] input_func_concat_DP5_0;
wire [31:0] input_func_concat_DP5_10;
wire [31:0] input_func_concat_DP5_11;
wire [31:0] input_func_concat_DP5_12;
wire [31:0] input_func_concat_DP5_13;
wire [31:0] input_func_concat_DP5_14;
wire [31:0] input_func_concat_DP5_15;
wire [31:0] input_func_concat_DP5_16;
wire [31:0] input_func_concat_DP5_17;
wire [31:0] input_func_concat_DP5_18;
wire [31:0] input_func_concat_DP5_19;
wire [31:0] input_func_concat_DP5_1;
wire [31:0] input_func_concat_DP5_20;
wire [31:0] input_func_concat_DP5_21;
wire [31:0] input_func_concat_DP5_22;
wire [31:0] input_func_concat_DP5_23;
wire [31:0] input_func_concat_DP5_24;
wire [31:0] input_func_concat_DP5_25;
wire [31:0] input_func_concat_DP5_26;
wire [31:0] input_func_concat_DP5_27;
wire [31:0] input_func_concat_DP5_28;
wire [31:0] input_func_concat_DP5_29;
wire [31:0] input_func_concat_DP5_2;
wire [31:0] input_func_concat_DP5_30;
wire [31:0] input_func_concat_DP5_31;
wire [31:0] input_func_concat_DP5_3;
wire [31:0] input_func_concat_DP5_4;
wire [31:0] input_func_concat_DP5_5;
wire [31:0] input_func_concat_DP5_6;
wire [31:0] input_func_concat_DP5_7;
wire [31:0] input_func_concat_DP5_8;
wire [31:0] input_func_concat_DP5_9;
wire [31:0] input_func_concat_DP6_0;
wire [31:0] input_func_concat_DP6_10;
wire [31:0] input_func_concat_DP6_11;
wire [31:0] input_func_concat_DP6_12;
wire [31:0] input_func_concat_DP6_13;
wire [31:0] input_func_concat_DP6_14;
wire [31:0] input_func_concat_DP6_15;
wire [31:0] input_func_concat_DP6_16;
wire [31:0] input_func_concat_DP6_17;
wire [31:0] input_func_concat_DP6_18;
wire [31:0] input_func_concat_DP6_19;
wire [31:0] input_func_concat_DP6_1;
wire [31:0] input_func_concat_DP6_20;
wire [31:0] input_func_concat_DP6_21;
wire [31:0] input_func_concat_DP6_22;
wire [31:0] input_func_concat_DP6_23;
wire [31:0] input_func_concat_DP6_24;
wire [31:0] input_func_concat_DP6_25;
wire [31:0] input_func_concat_DP6_26;
wire [31:0] input_func_concat_DP6_27;
wire [31:0] input_func_concat_DP6_2;
wire [31:0] input_func_concat_DP6_3;
wire [31:0] input_func_concat_DP6_4;
wire [31:0] input_func_concat_DP6_5;
wire [31:0] input_func_concat_DP6_6;
wire [31:0] input_func_concat_DP6_7;
wire [31:0] input_func_concat_DP6_8;
wire [31:0] input_func_concat_DP6_9;
wire [31:0] input_func_concat_DP7_0;
wire [31:0] input_func_concat_DP7_10;
wire [31:0] input_func_concat_DP7_11;
wire [31:0] input_func_concat_DP7_12;
wire [31:0] input_func_concat_DP7_13;
wire [31:0] input_func_concat_DP7_14;
wire [31:0] input_func_concat_DP7_15;
wire [31:0] input_func_concat_DP7_1;
wire [31:0] input_func_concat_DP7_2;
wire [31:0] input_func_concat_DP7_3;
wire [31:0] input_func_concat_DP7_4;
wire [31:0] input_func_concat_DP7_5;
wire [31:0] input_func_concat_DP7_6;
wire [31:0] input_func_concat_DP7_7;
wire [31:0] input_func_concat_DP7_8;
wire [31:0] input_func_concat_DP7_9;
wire [31:0] input_func_concat_MP0_0;
wire [31:0] input_func_concat_MP0_10;
wire [31:0] input_func_concat_MP0_11;
wire [31:0] input_func_concat_MP0_12;
wire [31:0] input_func_concat_MP0_13;
wire [31:0] input_func_concat_MP0_14;
wire [31:0] input_func_concat_MP0_15;
wire [31:0] input_func_concat_MP0_16;
wire [31:0] input_func_concat_MP0_17;
wire [31:0] input_func_concat_MP0_18;
wire [31:0] input_func_concat_MP0_19;
wire [31:0] input_func_concat_MP0_1;
wire [31:0] input_func_concat_MP0_20;
wire [31:0] input_func_concat_MP0_21;
wire [31:0] input_func_concat_MP0_22;
wire [31:0] input_func_concat_MP0_23;
wire [31:0] input_func_concat_MP0_24;
wire [31:0] input_func_concat_MP0_25;
wire [31:0] input_func_concat_MP0_26;
wire [31:0] input_func_concat_MP0_27;
wire [31:0] input_func_concat_MP0_28;
wire [31:0] input_func_concat_MP0_29;
wire [31:0] input_func_concat_MP0_2;
wire [31:0] input_func_concat_MP0_30;
wire [31:0] input_func_concat_MP0_31;
wire [31:0] input_func_concat_MP0_3;
wire [31:0] input_func_concat_MP0_4;
wire [31:0] input_func_concat_MP0_5;
wire [31:0] input_func_concat_MP0_6;
wire [31:0] input_func_concat_MP0_7;
wire [31:0] input_func_concat_MP0_8;
wire [31:0] input_func_concat_MP0_9;
wire [31:0] input_func_concat_MP1_0;
wire [31:0] input_func_concat_MP1_10;
wire [31:0] input_func_concat_MP1_11;
wire [31:0] input_func_concat_MP1_12;
wire [31:0] input_func_concat_MP1_13;
wire [31:0] input_func_concat_MP1_14;
wire [31:0] input_func_concat_MP1_15;
wire [31:0] input_func_concat_MP1_1;
wire [31:0] input_func_concat_MP1_2;
wire [31:0] input_func_concat_MP1_3;
wire [31:0] input_func_concat_MP1_4;
wire [31:0] input_func_concat_MP1_5;
wire [31:0] input_func_concat_MP1_6;
wire [31:0] input_func_concat_MP1_7;
wire [31:0] input_func_concat_MP1_8;
wire [31:0] input_func_concat_MP1_9;
wire [31:0] input_func_concat_MP2_0;
wire [31:0] input_func_concat_MP2_10;
wire [31:0] input_func_concat_MP2_11;
wire [31:0] input_func_concat_MP2_12;
wire [31:0] input_func_concat_MP2_13;
wire [31:0] input_func_concat_MP2_14;
wire [31:0] input_func_concat_MP2_15;
wire [31:0] input_func_concat_MP2_1;
wire [31:0] input_func_concat_MP2_2;
wire [31:0] input_func_concat_MP2_3;
wire [31:0] input_func_concat_MP2_4;
wire [31:0] input_func_concat_MP2_5;
wire [31:0] input_func_concat_MP2_6;
wire [31:0] input_func_concat_MP2_7;
wire [31:0] input_func_concat_MP2_8;
wire [31:0] input_func_concat_MP2_9;
assign input_func_concat_DP0_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4A_IN, `OUTPUTXBAR6_IN, `SPI8PICO_IN, `EPWM0A_IN, `TPIUCLK_IN, `CAN0TX_IN, 1'b0};
assign input_func_concat_DP0_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4B_IN, `OUTPUTXBAR7_IN, `SPI8POCI_IN, `EPWM0B_IN, `TPIUCTL_IN, `CAN0RX_IN, 1'b0};
assign input_func_concat_DP0_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5E_IN, `ADC0EXTMUXSEL0_IN, `SPI9CS1_IN, `EPWM5A_IN, `I2C2SDA_IN, `FSI0TXCLK_IN, 1'b0};
assign input_func_concat_DP0_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5F_IN, `ADC0EXTMUXSEL1_IN, `SPI9CS2_IN, `EPWM5B_IN, `I2C2SCL_IN, `FSI0TXD0_IN, 1'b0};
assign input_func_concat_DP0_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6A_IN, `nan_IN, `ADC0EXTMUXSEL2_IN, `SPI9CS3_IN, `EPWM6A_IN, `I2C3SDA_IN, `FSI0TXD1_IN, 1'b0};
assign input_func_concat_DP0_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6B_IN, `SPI9CS4_IN, `ADC0EXTMUXSEL3_IN, `FSI0TXCLK_IN, `EPWM6B_IN, `I2C3SCL_IN, `FSI0RXCLK_IN, 1'b0};
assign input_func_concat_DP0_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6C_IN, `SPI2CLK_IN, `MCPWM0A_IN, `FSI0TXD0_IN, `EPWM7A_IN, `RDC0PWM_N_IN, `FSI0RXD0_IN, 1'b0};
assign input_func_concat_DP0_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6D_IN, `SPI2PICO_IN, `MCPWM0B_IN, `FSI0TXD1_IN, `EPWM7B_IN, `RDC0PWM_P_IN, `FSI0RXD1_IN, 1'b0};
assign input_func_concat_DP0_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6E_IN, `SPI2POCI_IN, `MCPWM0C_IN, `FSI0RXCLK_IN, `EPWM8A_IN, `CLKOUT1_IN, `I2C0SDA_IN, 1'b0};
assign input_func_concat_DP0_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM6F_IN, `SPI2CS0_IN, `MCPWM0D_IN, `FSI0RXD0_IN, `EPWM8B_IN, `CLKOUT2_IN, `I2C0SCL_IN, 1'b0};
assign input_func_concat_DP0_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM7A_IN, `SPI2CS1_IN, `MCPWM0E_IN, `FSI0RXD1_IN, `EPWM9A_IN, `RDC1PWM_N_IN, `I2C1SDA_IN, 1'b0};
assign input_func_concat_DP0_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM7B_IN, `SPI2CS2_IN, `MCPWM0F_IN, `FSI1TXCLK_IN, `EPWM9B_IN, `RDC1PWM_P_IN, `I2C1SCL_IN, 1'b0};
assign input_func_concat_DP0_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4C_IN, `OUTPUTXBAR8_IN, `SPI8CS0_IN, `EPWM1A_IN, `TPIUDATA0_IN, `CAN1TX_IN, 1'b0};
assign input_func_concat_DP0_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS3_IN, `MCPWM1A_IN, `FSI1TXD0_IN, `EPWM10A_IN, `ADC2EXTMUXSEL0_IN, `LIN0TX_IN, 1'b0};
assign input_func_concat_DP0_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN4TX_IN, `MCPWM1B_IN, `FSI1TXD1_IN, `EPWM10B_IN, `ADC2EXTMUXSEL1_IN, `LIN0RX_IN, 1'b0};
assign input_func_concat_DP0_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN4RX_IN, `MCPWM1C_IN, `FSI1RXCLK_IN, `EPWM11A_IN, `ADC2EXTMUXSEL2_IN, `LIN1TX_IN, 1'b0};
assign input_func_concat_DP0_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN5TX_IN, `MCPWM1D_IN, `FSI1RXD0_IN, `EPWM11B_IN, `SPI7CS3_IN, `LIN1RX_IN, 1'b0};
assign input_func_concat_DP0_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN5RX_IN, `MCPWM1E_IN, `FSI1RXD1_IN, `EPWM12A_IN, `SPI7CLK_IN, `LIN2TX_IN, 1'b0};
assign input_func_concat_DP0_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS4_IN, `MCPWM1F_IN, `FSI2TXCLK_IN, `EPWM12B_IN, `SPI7PICO_IN, `LIN2RX_IN, 1'b0};
assign input_func_concat_DP0_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS5_IN, `OUTPUTXBAR0_IN, `FSI2TXD0_IN, `EPWM13A_IN, `SPI7POCI_IN, `LIN3TX_IN, 1'b0};
assign input_func_concat_DP0_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS5_IN, `OUTPUTXBAR1_IN, `FSI2TXD1_IN, `EPWM13B_IN, `SPI7CS0_IN, `LIN3RX_IN, 1'b0};
assign input_func_concat_DP0_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR2_IN, `FSI2RXCLK_IN, `EPWM14A_IN, `SPI7CS1_IN, `UART0TX_IN, 1'b0};
assign input_func_concat_DP0_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR3_IN, `FSI2RXD0_IN, `EPWM14B_IN, `SPI7CS2_IN, `UART0RX_IN, 1'b0};
assign input_func_concat_DP0_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4D_IN, `OUTPUTXBAR9_IN, `SPI8CS1_IN, `EPWM1B_IN, `TPIUDATA1_IN, `CAN1RX_IN, 1'b0};
assign input_func_concat_DP0_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR4_IN, `FSI2RXD1_IN, `EPWM15A_IN, `SPI5CLK_IN, `SENT0TXRX_IN, 1'b0};
assign input_func_concat_DP0_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR5_IN, `FSI3TXCLK_IN, `EPWM15B_IN, `SPI5PICO_IN, `SENT1TXRX_IN, 1'b0};
assign input_func_concat_DP0_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4E_IN, `OUTPUTXBAR10_IN, `SPI8CS2_IN, `EPWM2A_IN, `TPIUDATA2_IN, `CAN2TX_IN, 1'b0};
assign input_func_concat_DP0_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM4F_IN, `OUTPUTXBAR11_IN, `SPI8CS3_IN, `EPWM2B_IN, `TPIUDATA3_IN, `CAN2RX_IN, 1'b0};
assign input_func_concat_DP0_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5A_IN, `OUTPUTXBAR12_IN, `SPI9CLK_IN, `EPWM3A_IN, `ADC3EXTMUXSEL0_IN, `CAN3TX_IN, 1'b0};
assign input_func_concat_DP0_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5B_IN, `OUTPUTXBAR13_IN, `SPI9PICO_IN, `EPWM3B_IN, `ADC3EXTMUXSEL1_IN, `CAN3RX_IN, 1'b0};
assign input_func_concat_DP0_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5C_IN, `OUTPUTXBAR14_IN, `SPI9POCI_IN, `EPWM4A_IN, `ADC3EXTMUXSEL2_IN, `CAN4TX_IN, 1'b0};
assign input_func_concat_DP0_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM5D_IN, `OUTPUTXBAR15_IN, `SPI9CS0_IN, `EPWM4B_IN, `ADC3EXTMUXSEL3_IN, `CAN4RX_IN, 1'b0};
assign input_func_concat_DP1_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC0EXTMUXSEL0_IN, `FSI3RXCLK_IN, `SDFM0CLK_IN, `OUTPUTXBAR0_IN, `EPWM0A_IN, 1'b0};
assign input_func_concat_DP1_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC0EXTMUXSEL1_IN, `FSI3RXD0_IN, `SDFM0DATA_IN, `OUTPUTXBAR1_IN, `EPWM0B_IN, 1'b0};
assign input_func_concat_DP1_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SDFM5CLK_IN, `OUTPUTXBAR10_IN, `EPWM5A_IN, 1'b0};
assign input_func_concat_DP1_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SDFM5DATA_IN, `OUTPUTXBAR11_IN, `EPWM5B_IN, 1'b0};
assign input_func_concat_DP1_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SDFM6CLK_IN, `OUTPUTXBAR12_IN, `EPWM6A_IN, 1'b0};
assign input_func_concat_DP1_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN0TX_IN, `UART0TX_IN, `SDFM6DATA_IN, `OUTPUTXBAR13_IN, `EPWM6B_IN, 1'b0};
assign input_func_concat_DP1_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN0RX_IN, `UART0RX_IN, `SDFM7CLK_IN, `OUTPUTXBAR14_IN, `EPWM7A_IN, 1'b0};
assign input_func_concat_DP1_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN1TX_IN, `SPI8CLK_IN, `SDFM7DATA_IN, `OUTPUTXBAR15_IN, `EPWM7B_IN, 1'b0};
assign input_func_concat_DP1_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN1RX_IN, `SPI8PICO_IN, `SDFM8CLK_IN, `OUTPUTXBAR0_IN, `EPWM8A_IN, 1'b0};
assign input_func_concat_DP1_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN2TX_IN, `SPI8POCI_IN, `SDFM8DATA_IN, `OUTPUTXBAR1_IN, `EPWM8B_IN, 1'b0};
assign input_func_concat_DP1_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN2RX_IN, `SPI8CS0_IN, `SDFM9CLK_IN, `OUTPUTXBAR2_IN, `EPWM9A_IN, 1'b0};
assign input_func_concat_DP1_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN3TX_IN, `SPI8CS1_IN, `SDFM9DATA_IN, `OUTPUTXBAR3_IN, `EPWM9B_IN, 1'b0};
assign input_func_concat_DP1_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC0EXTMUXSEL2_IN, `FSI3RXD1_IN, `SDFM1CLK_IN, `OUTPUTXBAR2_IN, `EPWM1A_IN, 1'b0};
assign input_func_concat_DP1_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN3RX_IN, `SPI8CS2_IN, `SDFM10CLK_IN, `OUTPUTXBAR4_IN, `EPWM10A_IN, 1'b0};
assign input_func_concat_DP1_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS4_IN, `SPI8CS3_IN, `SDFM10DATA_IN, `OUTPUTXBAR5_IN, `EPWM10B_IN, 1'b0};
assign input_func_concat_DP1_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS5_IN, `SPI2CLK_IN, `SDFM11CLK_IN, `OUTPUTXBAR6_IN, `EPWM11A_IN, 1'b0};
assign input_func_concat_DP1_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2PICO_IN, `SDFM11DATA_IN, `OUTPUTXBAR7_IN, `EPWM11B_IN, 1'b0};
assign input_func_concat_DP1_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2POCI_IN, `ADC0EXTMUXSEL0_IN, `OUTPUTXBAR8_IN, `EPWM12A_IN, 1'b0};
assign input_func_concat_DP1_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS0_IN, `ADC0EXTMUXSEL1_IN, `OUTPUTXBAR9_IN, `EPWM12B_IN, 1'b0};
assign input_func_concat_DP1_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS1_IN, `ADC0EXTMUXSEL2_IN, `OUTPUTXBAR10_IN, `EPWM13A_IN, 1'b0};
assign input_func_concat_DP1_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS2_IN, `ADC0EXTMUXSEL3_IN, `OUTPUTXBAR11_IN, `EPWM13B_IN, 1'b0};
assign input_func_concat_DP1_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS3_IN, `ADC1EXTMUXSEL0_IN, `OUTPUTXBAR12_IN, `EPWM14A_IN, 1'b0};
assign input_func_concat_DP1_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CLK_IN, `ADC1EXTMUXSEL1_IN, `OUTPUTXBAR13_IN, `EPWM14B_IN, 1'b0};
assign input_func_concat_DP1_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC0EXTMUXSEL3_IN, `SPI8CS3_IN, `SDFM1DATA_IN, `OUTPUTXBAR3_IN, `EPWM1B_IN, 1'b0};
assign input_func_concat_DP1_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3PICO_IN, `ADC1EXTMUXSEL2_IN, `OUTPUTXBAR14_IN, `EPWM15A_IN, 1'b0};
assign input_func_concat_DP1_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3POCI_IN, `ADC1EXTMUXSEL3_IN, `OUTPUTXBAR15_IN, `EPWM15B_IN, 1'b0};
assign input_func_concat_DP1_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC2EXTMUXSEL0_IN, `SPI8CLK_IN, `SDFM2CLK_IN, `OUTPUTXBAR4_IN, `EPWM2A_IN, 1'b0};
assign input_func_concat_DP1_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC2EXTMUXSEL1_IN, `SPI8PICO_IN, `SDFM2DATA_IN, `OUTPUTXBAR5_IN, `EPWM2B_IN, 1'b0};
assign input_func_concat_DP1_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC2EXTMUXSEL2_IN, `SPI8POCI_IN, `SDFM3CLK_IN, `OUTPUTXBAR6_IN, `EPWM3A_IN, 1'b0};
assign input_func_concat_DP1_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC2EXTMUXSEL3_IN, `SPI8CS0_IN, `SDFM3DATA_IN, `OUTPUTXBAR7_IN, `EPWM3B_IN, 1'b0};
assign input_func_concat_DP1_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI8CS1_IN, `SDFM4CLK_IN, `OUTPUTXBAR8_IN, `EPWM4A_IN, 1'b0};
assign input_func_concat_DP1_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI8CS2_IN, `SDFM4DATA_IN, `OUTPUTXBAR9_IN, `EPWM4B_IN, 1'b0};
assign input_func_concat_DP2_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS0_IN, `ADC2EXTMUXSEL0_IN, `CLKOUT1_IN, `EPWM16A_IN, 1'b0};
assign input_func_concat_DP2_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS1_IN, `ADC2EXTMUXSEL1_IN, `ADC4EXTMUXSEL0_IN, `EPWM16B_IN, 1'b0};
assign input_func_concat_DP2_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS3_IN, `ADC4EXTMUXSEL2_IN, `CLKOUT2_IN, `EPWM21A_IN, 1'b0};
assign input_func_concat_DP2_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CLK_IN, `ADC4EXTMUXSEL3_IN, `nan_IN, `EPWM21B_IN, 1'b0};
assign input_func_concat_DP2_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1TXCLK_IN, `nan_IN, `SPI5PICO_IN, `ADC5EXTMUXSEL0_IN, `MCASP0EXTREFCLK_IN, `EPWM22A_IN, 1'b0};
assign input_func_concat_DP2_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1TXD0_IN, `I2C0SDA_IN, `SPI5POCI_IN, `ADC5EXTMUXSEL1_IN, `MCASP0ACLKX_IN, `EPWM22B_IN, 1'b0};
assign input_func_concat_DP2_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1TXD1_IN, `I2C0SCL_IN, `SPI5CS0_IN, `ADC5EXTMUXSEL2_IN, `MCASP0AFSX_IN, `EPWM23A_IN, 1'b0};
assign input_func_concat_DP2_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1RXCLK_IN, `I2C1SDA_IN, `SPI5CS1_IN, `ADC5EXTMUXSEL3_IN, `MCASP0ACLKR_IN, `EPWM23B_IN, 1'b0};
assign input_func_concat_DP2_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1RXD0_IN, `I2C1SCL_IN, `SPI5CS2_IN, `ADC6EXTMUXSEL0_IN, `MCASP0AFSR_IN, `EPWM24A_IN, 1'b0};
assign input_func_concat_DP2_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI1RXD1_IN, `I2C2SDA_IN, `SPI5CS3_IN, `ADC6EXTMUXSEL1_IN, `MCASP0AXR0_IN, `EPWM24B_IN, 1'b0};
assign input_func_concat_DP2_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI2TXCLK_IN, `I2C2SCL_IN, `SPI6CLK_IN, `ADC6EXTMUXSEL2_IN, `MCASP0AXR1_IN, `EPWM25A_IN, 1'b0};
assign input_func_concat_DP2_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI2TXD0_IN, `I2C3SDA_IN, `SPI6PICO_IN, `ADC6EXTMUXSEL3_IN, `MCASP0AXR2_IN, `EPWM25B_IN, 1'b0};
assign input_func_concat_DP2_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS2_IN, `ADC2EXTMUXSEL2_IN, `ADC4EXTMUXSEL1_IN, `EPWM17A_IN, 1'b0};
assign input_func_concat_DP2_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `FSI2TXD1_IN, `I2C3SCL_IN, `SPI6POCI_IN, `ADC7EXTMUXSEL0_IN, `MCASP0AXR3_IN, `EPWM26A_IN, 1'b0};
assign input_func_concat_DP2_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2A_IN, `SPI8CS4_IN, `SPI6CS0_IN, `ADC7EXTMUXSEL1_IN, `CAN6TX_IN, `EPWM26B_IN, 1'b0};
assign input_func_concat_DP2_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2B_IN, `SPI8CS5_IN, `SPI6CS1_IN, `ADC7EXTMUXSEL2_IN, `CAN6RX_IN, `EPWM27A_IN, 1'b0};
assign input_func_concat_DP2_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2C_IN, `SPI3CS4_IN, `SPI6CS2_IN, `ADC7EXTMUXSEL3_IN, `CAN7TX_IN, `EPWM27B_IN, 1'b0};
assign input_func_concat_DP2_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2D_IN, `SPI3CS5_IN, `SPI6CS3_IN, `ADCSOC0_IN, `CAN7RX_IN, `EPWM28A_IN, 1'b0};
assign input_func_concat_DP2_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2E_IN, `LIN6TX_IN, `SPI7CLK_IN, `ADCSOC1_IN, `CAN8TX_IN, `EPWM28B_IN, 1'b0};
assign input_func_concat_DP2_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM2F_IN, `LIN6RX_IN, `SPI7PICO_IN, `SPI6CLK_IN, `CAN8RX_IN, `EPWM29A_IN, 1'b0};
assign input_func_concat_DP2_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3A_IN, `LIN7TX_IN, `SPI7POCI_IN, `SPI6PICO_IN, `CAN9TX_IN, `EPWM29B_IN, 1'b0};
assign input_func_concat_DP2_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3B_IN, `LIN7RX_IN, `SPI7CS0_IN, `SPI6POCI_IN, `CAN9RX_IN, `EPWM30A_IN, 1'b0};
assign input_func_concat_DP2_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3C_IN, `SDFM7CLK_IN, `SPI7CS1_IN, `SPI6CS0_IN, `CAN10TX_IN, `EPWM30B_IN, 1'b0};
assign input_func_concat_DP2_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS3_IN, `ADC2EXTMUXSEL3_IN, `ADC4EXTMUXSEL2_IN, `EPWM17B_IN, 1'b0};
assign input_func_concat_DP2_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3D_IN, `SDFM7DATA_IN, `SPI7CS2_IN, `SPI6CS1_IN, `CAN10RX_IN, `EPWM31A_IN, 1'b0};
assign input_func_concat_DP2_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3E_IN, `SDFM0CLK_IN, `SPI7CS3_IN, `SPI6CS2_IN, `CAN11TX_IN, `EPWM31B_IN, 1'b0};
assign input_func_concat_DP2_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CLK_IN, `ADC3EXTMUXSEL0_IN, `ADC4EXTMUXSEL3_IN, `EPWM18A_IN, 1'b0};
assign input_func_concat_DP2_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4PICO_IN, `ADC3EXTMUXSEL1_IN, `ADC5EXTMUXSEL0_IN, `EPWM18B_IN, 1'b0};
assign input_func_concat_DP2_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4POCI_IN, `ADC3EXTMUXSEL2_IN, `ADC5EXTMUXSEL1_IN, `EPWM19A_IN, 1'b0};
assign input_func_concat_DP2_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS0_IN, `ADC3EXTMUXSEL3_IN, `ADC5EXTMUXSEL2_IN, `EPWM19B_IN, 1'b0};
assign input_func_concat_DP2_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS1_IN, `ADC4EXTMUXSEL0_IN, `ADC5EXTMUXSEL3_IN, `EPWM20A_IN, 1'b0};
assign input_func_concat_DP2_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS2_IN, `ADC4EXTMUXSEL1_IN, `CLKOUT1_IN, `EPWM20B_IN, 1'b0};
assign input_func_concat_DP3_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM3F_IN, `SDFM0DATA_IN, `SPI8CLK_IN, `SPI6CS3_IN, `CAN11RX_IN, `EPWMSYNCO_IN, 1'b0};
assign input_func_concat_DP3_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC3EXTMUXSEL0_IN, `SPI4CLK_IN, `FSI3TXD0_IN, `EPWM16A_IN, `SPI5POCI_IN, `SENT2TXRX_IN, 1'b0};
assign input_func_concat_DP3_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_TX_IN, `SPI5POCI_IN, `FSI4RXD0_IN, `EPWM20B_IN, `SPI4POCI_IN, `MIBSPI0CS3_IN, 1'b0};
assign input_func_concat_DP3_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_RX_IN, `SPI5CS0_IN, `FSI4RXD1_IN, `EPWM21A_IN, `SPI3CS5_IN, `MIBSPI1CLK_IN, 1'b0};
assign input_func_concat_DP3_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_TX_IN, `SPI5CS1_IN, `FSI5TXCLK_IN, `EPWM21B_IN, `MCPWM10A_IN, `MIBSPI1PICO_IN, 1'b0};
assign input_func_concat_DP3_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_RX_IN, `SPI5CS2_IN, `FSI5TXD0_IN, `EPWM22A_IN, `MCPWM10B_IN, `MIBSPI1POCI_IN, 1'b0};
assign input_func_concat_DP3_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS4_IN, `SPI5CS3_IN, `FSI5TXD1_IN, `EPWM22B_IN, `ADC2EXTMUXSEL3_IN, `MIBSPI1CS0_IN, 1'b0};
assign input_func_concat_DP3_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS5_IN, `SPI6CLK_IN, `FSI5RXCLK_IN, `EPWM23A_IN, `SPI4CS0_IN, `MIBSPI1CS1_IN, 1'b0};
assign input_func_concat_DP3_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS6_IN, `SPI6PICO_IN, `FSI5RXD0_IN, `EPWM23B_IN, `SPI4CS1_IN, `MIBSPI1CS2_IN, 1'b0};
assign input_func_concat_DP3_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS7_IN, `SPI6POCI_IN, `FSI5RXD1_IN, `EPWM24A_IN, `SPI4CS2_IN, `MCPWM0A_IN, 1'b0};
assign input_func_concat_DP3_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS8_IN, `SPI6CS0_IN, `MCPWM7E_IN, `EPWM24B_IN, `SPI4CS3_IN, `MCPWM0B_IN, 1'b0};
assign input_func_concat_DP3_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS9_IN, `SPI6CS1_IN, `MCPWM7F_IN, `EPWM25A_IN, `ADC1EXTMUXSEL0_IN, `MCPWM0C_IN, 1'b0};
assign input_func_concat_DP3_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC3EXTMUXSEL1_IN, `SPI4PICO_IN, `FSI3TXD1_IN, `EPWM16B_IN, `SPI5CS0_IN, `SENT3TXRX_IN, 1'b0};
assign input_func_concat_DP3_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS10_IN, `SPI6CS2_IN, `MCPWM8A_IN, `EPWM25B_IN, `ADC1EXTMUXSEL1_IN, `MCPWM0D_IN, 1'b0};
assign input_func_concat_DP3_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS11_IN, `SPI6CS3_IN, `MCPWM8B_IN, `EPWM26A_IN, `ADC1EXTMUXSEL2_IN, `MCPWM0E_IN, 1'b0};
assign input_func_concat_DP3_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CLK_IN, `EPWM31B_IN, `MCPWM8C_IN, `EPWM26B_IN, `ADC1EXTMUXSEL3_IN, `MCPWM0F_IN, 1'b0};
assign input_func_concat_DP3_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3PICO_IN, `EPWM31A_IN, `MCPWM8D_IN, `EPWM27A_IN, `FSI5TXCLK_IN, `MCPWM1A_IN, 1'b0};
assign input_func_concat_DP3_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3POCI_IN, `EPWM30B_IN, `MCPWM8E_IN, `EPWM27B_IN, `FSI5TXD0_IN, `MCPWM1B_IN, 1'b0};
assign input_func_concat_DP3_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS0_IN, `EPWM30A_IN, `MCPWM8F_IN, `EPWM28A_IN, `FSI5TXD1_IN, `MCPWM1C_IN, 1'b0};
assign input_func_concat_DP3_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS1_IN, `EPWM29B_IN, `MCPWM9A_IN, `EPWM28B_IN, `FSI5RXCLK_IN, `MCPWM1D_IN, 1'b0};
assign input_func_concat_DP3_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS2_IN, `EPWM29A_IN, `MCPWM9B_IN, `EPWM29A_IN, `FSI5RXD0_IN, `MCPWM1E_IN, 1'b0};
assign input_func_concat_DP3_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI3CS3_IN, `EPWM28B_IN, `MCPWM9C_IN, `EPWM29B_IN, `FSI5RXD1_IN, `MCPWM1F_IN, 1'b0};
assign input_func_concat_DP3_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM28A_IN, `MCPWM9D_IN, `I2C0SDA_IN, `SPI8CLK_IN, `MIBSPI1CS3_IN, 1'b0};
assign input_func_concat_DP3_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC3EXTMUXSEL2_IN, `SPI4POCI_IN, `FSI3RXCLK_IN, `EPWM17A_IN, `SPI5CS1_IN, `SENT4TXRX_IN, 1'b0};
assign input_func_concat_DP3_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM27B_IN, `MCPWM9E_IN, `I2C0SCL_IN, `SPI8PICO_IN, `PSI5_0_TX_IN, 1'b0};
assign input_func_concat_DP3_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM27A_IN, `MCPWM9F_IN, `I2C1SDA_IN, `SPI8POCI_IN, `PSI5_0_RX_IN, 1'b0};
assign input_func_concat_DP3_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC3EXTMUXSEL3_IN, `SPI4CS0_IN, `FSI3RXD0_IN, `EPWM17B_IN, `SPI5CS2_IN, `MIBSPI0CLK_IN, 1'b0};
assign input_func_concat_DP3_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS1_IN, `FSI3RXD1_IN, `EPWM18A_IN, `SPI5CS3_IN, `MIBSPI0PICO_IN, 1'b0};
assign input_func_concat_DP3_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS2_IN, `FSI4TXCLK_IN, `EPWM18B_IN, `SPI3CS4_IN, `MIBSPI0POCI_IN, 1'b0};
assign input_func_concat_DP3_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS3_IN, `FSI4TXD0_IN, `EPWM19A_IN, `EXTCLK_IN, `MIBSPI0CS0_IN, 1'b0};
assign input_func_concat_DP3_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CLK_IN, `FSI4TXD1_IN, `EPWM19B_IN, `SPI4CLK_IN, `MIBSPI0CS1_IN, 1'b0};
assign input_func_concat_DP3_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5PICO_IN, `FSI4RXCLK_IN, `EPWM20A_IN, `SPI4PICO_IN, `MIBSPI0CS2_IN, 1'b0};
assign input_func_concat_DP4_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM26B_IN, `MCPWM10A_IN, `I2C1SCL_IN, `SPI8CS0_IN, `PSI5_1_TX_IN, 1'b0};
assign input_func_concat_DP4_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM26A_IN, `MCPWM10B_IN, `I2C2SDA_IN, `SPI8CS1_IN, `PSI5_1_RX_IN, 1'b0};
assign input_func_concat_DP4_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC7EXTMUXSEL0_IN, `MIBSPI0POCI_IN, `EPWM21B_IN, `MCASP0AFSR_IN, `MCPWM6E_IN, `PSI5_1_TX_IN, `RGMII1TXD3_IN, 1'b0};
assign input_func_concat_DP4_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC7EXTMUXSEL1_IN, `MIBSPI0CS0_IN, `EPWM21A_IN, `MCASP0AXR0_IN, `MCPWM6F_IN, `PSI5_1_RX_IN, `RGMII1TXCTL_IN, 1'b0};
assign input_func_concat_DP4_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC7EXTMUXSEL2_IN, `MIBSPI0CS1_IN, `EPWM20B_IN, `MCASP0AXR1_IN, `MCPWM7A_IN, `FSI4TXCLK_IN, `RGMII1RXCLK_IN, 1'b0};
assign input_func_concat_DP4_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC7EXTMUXSEL3_IN, `MIBSPI0CS2_IN, `EPWM20A_IN, `MCASP0AXR2_IN, `MCPWM7B_IN, `FSI4TXD0_IN, `RGMII1RXD0_IN, 1'b0};
assign input_func_concat_DP4_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS3_IN, `EPWM19B_IN, `MCASP0AXR3_IN, `MCPWM7C_IN, `FSI4TXD1_IN, `RGMII1RXD1_IN, 1'b0};
assign input_func_concat_DP4_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS4_IN, `SENT0TXRX_IN, `EPWM19A_IN, `MCPWM9D_IN, `MCPWM7D_IN, `FSI4RXCLK_IN, `RGMII1RXD2_IN, 1'b0};
assign input_func_concat_DP4_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS5_IN, `SENT1TXRX_IN, `EPWM18B_IN, `MCPWM9E_IN, `MCPWM7E_IN, `FSI4RXD0_IN, `RGMII1RXD3_IN, 1'b0};
assign input_func_concat_DP4_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS6_IN, `SENT2TXRX_IN, `EPWM18A_IN, `MCPWM9F_IN, `MCPWM7F_IN, `FSI4RXD1_IN, `RGMII1RXCTL_IN, 1'b0};
assign input_func_concat_DP4_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM17B_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS4_IN, 1'b0};
assign input_func_concat_DP4_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM17A_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS5_IN, 1'b0};
assign input_func_concat_DP4_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM25B_IN, `MCPWM10C_IN, `I2C2SCL_IN, `SPI8CS2_IN, `SPI3CLK_IN, 1'b0};
assign input_func_concat_DP4_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS7_IN, `MIBSPI1CLK_IN, `EPWM16B_IN, `MCASP0EXTREFCLK_IN, `EPWM30A_IN, `RDC0PWM_N_IN, `XSPI0CLK_IN, 1'b0};
assign input_func_concat_DP4_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS8_IN, `MIBSPI1PICO_IN, `EPWM16A_IN, `MCASP0ACLKX_IN, `EPWM30B_IN, `RDC0PWM_P_IN, `XSPI0CS0_IN, 1'b0};
assign input_func_concat_DP4_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS9_IN, `MIBSPI1POCI_IN, `EPWM15B_IN, `MCASP0AFSX_IN, `EPWM31A_IN, `RDC1PWM_N_IN, `XSPI0CS1_IN, 1'b0};
assign input_func_concat_DP4_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS10_IN, `MIBSPI1CS0_IN, `EPWM15A_IN, `MCASP0ACLKR_IN, `EPWM31B_IN, `RDC1PWM_P_IN, `XSPI0DS0_IN, 1'b0};
assign input_func_concat_DP4_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS11_IN, `MIBSPI1CS1_IN, `EPWM14B_IN, `MCASP0AFSR_IN, `EPWMSYNCO_IN, `LIN4TX_IN, `XSPI0DS1_IN, 1'b0};
assign input_func_concat_DP4_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS2_IN, `EPWM14A_IN, `MCASP0AXR0_IN, `SPI2CS4_IN, `LIN4RX_IN, `XSPI0DS2_IN, 1'b0};
assign input_func_concat_DP4_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS3_IN, `EPWM13B_IN, `MCASP0AXR1_IN, `MCPWM10A_IN, `LIN5TX_IN, `XSPI0DS3_IN, 1'b0};
assign input_func_concat_DP4_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS5_IN, `EPWM13A_IN, `MCASP0AXR2_IN, `MCPWM10B_IN, `LIN5RX_IN, `XSPI0DS4_IN, 1'b0};
assign input_func_concat_DP4_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN0TX_IN, `EPWM12B_IN, `MCASP0AXR3_IN, `MCPWM10C_IN, `LIN6TX_IN, `XSPI0DS5_IN, 1'b0};
assign input_func_concat_DP4_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN0RX_IN, `EPWM12A_IN, `MSC0CLK_IN, `MCPWM10D_IN, `LIN6RX_IN, `XSPI0DS6_IN, 1'b0};
assign input_func_concat_DP4_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM25A_IN, `MCPWM10D_IN, `I2C3SDA_IN, `SPI8CS3_IN, `SPI3PICO_IN, 1'b0};
assign input_func_concat_DP4_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CLK_IN, `CAN1TX_IN, `EPWM11B_IN, `MSC0SI_IN, `MCPWM10E_IN, `SENT5TXRX_IN, `XSPI0DS7_IN, 1'b0};
assign input_func_concat_DP4_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4PICO_IN, `CAN1RX_IN, `EPWM11A_IN, `MSC0SO_IN, `MCPWM10F_IN, `EXTCLK_IN, `XSPI0DQS_IN, 1'b0};
assign input_func_concat_DP4_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS4_IN, `EPWM24B_IN, `MCPWM10E_IN, `I2C3SCL_IN, `nan_IN, `SPI3POCI_IN, 1'b0};
assign input_func_concat_DP4_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI2CS5_IN, `EPWM24A_IN, `MCPWM10F_IN, `nan_IN, `SPI3CS1_IN, `SPI3CS0_IN, 1'b0};
assign input_func_concat_DP4_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC6EXTMUXSEL0_IN, `UART1TX_IN, `EPWM23B_IN, `MCASP0EXTREFCLK_IN, `MCPWM6A_IN, `SPI3CS2_IN, `RGMII1TXCLK_IN, 1'b0};
assign input_func_concat_DP4_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC6EXTMUXSEL1_IN, `UART1RX_IN, `EPWM23A_IN, `MCASP0ACLKX_IN, `MCPWM6B_IN, `SPI3CS3_IN, `RGMII1TXD0_IN, 1'b0};
assign input_func_concat_DP4_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC6EXTMUXSEL2_IN, `MIBSPI0CLK_IN, `EPWM22B_IN, `MCASP0AFSX_IN, `MCPWM6C_IN, `PSI5_0_TX_IN, `RGMII1TXD1_IN, 1'b0};
assign input_func_concat_DP4_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `ADC6EXTMUXSEL3_IN, `MIBSPI0PICO_IN, `EPWM22A_IN, `MCASP0ACLKR_IN, `MCPWM6D_IN, `PSI5_0_RX_IN, `RGMII1TXD2_IN, 1'b0};
assign input_func_concat_DP5_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4POCI_IN, `PSI5_0_TX_IN, `EPWM10B_IN, `MSC0CS0_IN, `MCPWM7C_IN, `MIBSPI0CS2_IN, `GMII_MDC_IN, 1'b0};
assign input_func_concat_DP5_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS0_IN, `PSI5_0_RX_IN, `EPWM10A_IN, `MSC0CS1_IN, `MCPWM7D_IN, `MIBSPI0CS3_IN, `GMII_MDIO_IN, 1'b0};
assign input_func_concat_DP5_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS0_IN, `EPWM5B_IN, `SPI2CS0_IN, `MCPWM3C_IN, `MIBSPI0PICO_IN, `RGMII0RXD1_IN, 1'b0};
assign input_func_concat_DP5_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS1_IN, `EPWM5A_IN, `SPI2CS1_IN, `MCPWM3D_IN, `MIBSPI0POCI_IN, `RGMII0RXD2_IN, 1'b0};
assign input_func_concat_DP5_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS2_IN, `EPWM4B_IN, `SPI2CS2_IN, `MCPWM3E_IN, `MIBSPI0CS0_IN, `RGMII0RXD3_IN, 1'b0};
assign input_func_concat_DP5_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS3_IN, `EPWM4A_IN, `SPI2CS3_IN, `MCPWM3F_IN, `MIBSPI0CS1_IN, `RGMII0RXCTL_IN, 1'b0};
assign input_func_concat_DP5_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CLK_IN, `EPWM3B_IN, `MCPWM0A_IN, `RDC0PWM_N_IN, `CAN0TX_IN, `TPIUCLK_IN, 1'b0};
assign input_func_concat_DP5_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7PICO_IN, `EPWM3A_IN, `MCPWM0B_IN, `RDC0PWM_P_IN, `CAN0RX_IN, `TPIUCTL_IN, 1'b0};
assign input_func_concat_DP5_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7POCI_IN, `EPWM2B_IN, `MCPWM0C_IN, `RDC1PWM_N_IN, `CAN1TX_IN, `TPIUDATA0_IN, 1'b0};
assign input_func_concat_DP5_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS0_IN, `EPWM2A_IN, `MCPWM0D_IN, `RDC1PWM_P_IN, `CAN1RX_IN, `TPIUDATA1_IN, 1'b0};
assign input_func_concat_DP5_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS1_IN, `EPWM1B_IN, `MCPWM0E_IN, `nan_IN, `CAN2TX_IN, `TPIUDATA2_IN, 1'b0};
assign input_func_concat_DP5_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS2_IN, `EPWM1A_IN, `MCPWM0F_IN, `nan_IN, `CAN2RX_IN, `TPIUDATA3_IN, 1'b0};
assign input_func_concat_DP5_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS1_IN, `PSI5_1_TX_IN, `EPWM9B_IN, `MSC0CS2_IN, `MCPWM2A_IN, `SPI9CLK_IN, `RGMII0TXCLK_IN, 1'b0};
assign input_func_concat_DP5_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS3_IN, `EPWM0B_IN, `MCPWM1A_IN, `ADC6EXTMUXSEL0_IN, `CAN3TX_IN, `SPI2CLK_IN, 1'b0};
assign input_func_concat_DP5_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_TX_IN, `EPWM0A_IN, `MCPWM1B_IN, `ADC6EXTMUXSEL1_IN, `CAN3RX_IN, `SPI2PICO_IN, 1'b0};
assign input_func_concat_DP5_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_RX_IN, `EPWM0A_IN, `MCPWM1C_IN, `ADC7EXTMUXSEL0_IN, `CAN4TX_IN, `SPI2POCI_IN, 1'b0};
assign input_func_concat_DP5_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS1_IN, `PSI5_2_TX_IN, `MCPWM1D_IN, `ADC7EXTMUXSEL1_IN, `CAN4RX_IN, `SPI2CS0_IN, 1'b0};
assign input_func_concat_DP5_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS2_IN, `PSI5_2_RX_IN, `MCPWM1E_IN, `ADC7EXTMUXSEL2_IN, `SPI2CS1_IN, `CAN5TX_IN, 1'b0};
assign input_func_concat_DP5_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS3_IN, `nan_IN, `MCPWM1F_IN, `ADC7EXTMUXSEL3_IN, `SPI2CS2_IN, `CAN5RX_IN, 1'b0};
assign input_func_concat_DP5_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM24A_IN, `MIBSPI1CLK_IN, `MCPWM2A_IN, `MCPWM4A_IN, `SPI2CS3_IN, `RGMII2TXCLK_IN, 1'b0};
assign input_func_concat_DP5_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_TX_IN, `EPWM24B_IN, `MIBSPI1PICO_IN, `MCPWM2B_IN, `MCPWM4B_IN, `FSI1TXCLK_IN, `RGMII2TXD0_IN, 1'b0};
assign input_func_concat_DP5_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_RX_IN, `EPWM25A_IN, `MIBSPI1POCI_IN, `MCPWM2C_IN, `MCPWM4C_IN, `FSI1TXD0_IN, `RGMII2TXD1_IN, 1'b0};
assign input_func_concat_DP5_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_TX_IN, `EPWM25B_IN, `MIBSPI1CS0_IN, `MCPWM2D_IN, `MCPWM4D_IN, `FSI1TXD1_IN, `RGMII2TXD2_IN, 1'b0};
assign input_func_concat_DP5_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS2_IN, `PSI5_1_RX_IN, `EPWM9A_IN, `MSC0CS3_IN, `MCPWM2B_IN, `SPI9PICO_IN, `RGMII0TXD0_IN, 1'b0};
assign input_func_concat_DP5_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_RX_IN, `EPWM26A_IN, `MIBSPI1CS1_IN, `MCPWM2E_IN, `MCPWM4E_IN, `FSI1RXCLK_IN, `RGMII2TXD3_IN, 1'b0};
assign input_func_concat_DP5_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_TX_IN, `SPI9CLK_IN, `EPWM26B_IN, `MIBSPI1CS2_IN, `MCPWM2F_IN, `MCPWM4F_IN, `FSI1RXD0_IN, `RGMII2TXCTL_IN, 1'b0};
assign input_func_concat_DP5_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS3_IN, `SENT3TXRX_IN, `EPWM8B_IN, `LIN7TX_IN, `MCPWM2C_IN, `SPI9POCI_IN, `RGMII0TXD1_IN, 1'b0};
assign input_func_concat_DP5_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SENT4TXRX_IN, `EPWM8A_IN, `LIN7RX_IN, `MCPWM2D_IN, `SPI9CS0_IN, `RGMII0TXD2_IN, 1'b0};
assign input_func_concat_DP5_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SENT5TXRX_IN, `EPWM7B_IN, `MIBSPI1CS3_IN, `MCPWM2E_IN, `SPI9CS1_IN, `RGMII0TXD3_IN, 1'b0};
assign input_func_concat_DP5_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CLK_IN, `EPWM7A_IN, `SPI2CLK_IN, `MCPWM2F_IN, `SPI9CS2_IN, `RGMII0TXCTL_IN, 1'b0};
assign input_func_concat_DP5_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6PICO_IN, `EPWM6B_IN, `SPI2PICO_IN, `MCPWM3A_IN, `SPI9CS3_IN, `RGMII0RXCLK_IN, 1'b0};
assign input_func_concat_DP5_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6POCI_IN, `EPWM6A_IN, `SPI2POCI_IN, `MCPWM3B_IN, `MIBSPI0CLK_IN, `RGMII0RXD0_IN, 1'b0};
assign input_func_concat_DP6_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_2_RX_IN, `SPI9PICO_IN, `SPI5CLK_IN, `MIBSPI1CS3_IN, `MCPWM3A_IN, `MCPWM5A_IN, `FSI1RXD1_IN, `RGMII2RXCLK_IN, 1'b0};
assign input_func_concat_DP6_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_TX_IN, `SPI9POCI_IN, `SPI5PICO_IN, `nan_IN, `MCPWM3B_IN, `MCPWM5B_IN, `FSI2TXCLK_IN, `RGMII2RXD0_IN, 1'b0};
assign input_func_concat_DP6_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR6_IN, `EPWM3A_IN, `MSC1CS1_IN, `MCPWM4E_IN, `MCPWM8E_IN, `FSI3TXD0_IN, `MMC0DATA2_IN, 1'b0};
assign input_func_concat_DP6_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR7_IN, `EPWM3B_IN, `MSC1CS2_IN, `MCPWM4F_IN, `MCPWM8F_IN, `FSI3TXD1_IN, `MMC0DATA3_IN, 1'b0};
assign input_func_concat_DP6_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR8_IN, `EPWM24A_IN, `MSC1CS3_IN, `MCPWM5A_IN, `MSC1CLK_IN, `CAN5TX_IN, `MMC0CD_IN, 1'b0};
assign input_func_concat_DP6_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR9_IN, `EPWM24B_IN, `CLKOUT2_IN, `MCPWM5B_IN, `MSC1SI_IN, `CAN5RX_IN, `MMC0WP_IN, 1'b0};
assign input_func_concat_DP6_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR10_IN, `EPWM25A_IN, `ADC4EXTMUXSEL0_IN, `MCPWM5C_IN, `MSC1SO_IN, `MSC0CLK_IN, `T1S0TX_IN, 1'b0};
assign input_func_concat_DP6_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR11_IN, `EPWM25B_IN, `ADC4EXTMUXSEL1_IN, `MCPWM5D_IN, `MSC1CS0_IN, `MSC0SI_IN, `T1S0RX_IN, 1'b0};
assign input_func_concat_DP6_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR12_IN, `EPWM26A_IN, `ADC4EXTMUXSEL2_IN, `MCPWM5E_IN, `MSC1CS1_IN, `MSC0SO_IN, `T1S0ED_IN, 1'b0};
assign input_func_concat_DP6_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR13_IN, `EPWM26B_IN, `ADC4EXTMUXSEL3_IN, `MCPWM5F_IN, `MSC1CS2_IN, `MSC0CS0_IN, `T1S1TX_IN, 1'b0};
assign input_func_concat_DP6_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS4_IN, `CAN2TX_IN, `CLKOUT2_IN, `MCPWM6A_IN, `MSC1CS3_IN, `MSC0CS1_IN, `T1S1RX_IN, 1'b0};
assign input_func_concat_DP6_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS5_IN, `CAN2RX_IN, `SPI3CLK_IN, `MCPWM6B_IN, `CLKOUT1_IN, `MSC0CS2_IN, `T1S1ED_IN, 1'b0};
assign input_func_concat_DP6_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `PSI5_3_RX_IN, `SPI9CS0_IN, `SPI5POCI_IN, `ADC5EXTMUXSEL0_IN, `MCPWM3C_IN, `MCPWM5C_IN, `FSI2TXD0_IN, `RGMII2RXD1_IN, 1'b0};
assign input_func_concat_DP6_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS6_IN, `CAN3TX_IN, `SPI3PICO_IN, `MCPWM6C_IN, `MCPWM9A_IN, `MSC1CLK_IN, `T1S2TX_IN, 1'b0};
assign input_func_concat_DP6_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS7_IN, `CAN3RX_IN, `SPI3POCI_IN, `MCPWM6D_IN, `MCPWM9B_IN, `MSC1SI_IN, `T1S2RX_IN, 1'b0};
assign input_func_concat_DP6_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS8_IN, `CAN4TX_IN, `SPI3CS0_IN, `MCPWM6E_IN, `MCPWM9C_IN, `MSC1SO_IN, `T1S2ED_IN, 1'b0};
assign input_func_concat_DP6_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS9_IN, `CAN4RX_IN, `SPI3CS1_IN, `MCPWM6F_IN, `MCPWM9D_IN, `MSC1CS0_IN, `T1S3TX_IN, 1'b0};
assign input_func_concat_DP6_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS10_IN, `CAN5TX_IN, `SPI3CS2_IN, `MCPWM7A_IN, `MCPWM9E_IN, `MSC1CS1_IN, `T1S3RX_IN, 1'b0};
assign input_func_concat_DP6_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS11_IN, `CAN5RX_IN, `SPI3CS3_IN, `MCPWM7B_IN, `MCPWM9F_IN, `MSC0CS3_IN, `T1S3ED_IN, 1'b0};
assign input_func_concat_DP6_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM7C_IN, `ADC6EXTMUXSEL2_IN, `MSC1CS2_IN, `T1SMDC_IN, 1'b0};
assign input_func_concat_DP6_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM7D_IN, `ADC6EXTMUXSEL3_IN, `MSC1CS3_IN, `T1SMDIO_IN, 1'b0};
assign input_func_concat_DP6_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS1_IN, `SPI5CS0_IN, `ADC5EXTMUXSEL1_IN, `MCPWM3D_IN, `MCPWM5D_IN, `FSI2TXD1_IN, `RGMII2RXD2_IN, 1'b0};
assign input_func_concat_DP6_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS2_IN, `nan_IN, `ADC5EXTMUXSEL2_IN, `MCPWM3E_IN, `MCPWM5E_IN, `ADCSOC0_IN, `RGMII2RXD3_IN, 1'b0};
assign input_func_concat_DP6_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS3_IN, `nan_IN, `ADC5EXTMUXSEL3_IN, `MCPWM3F_IN, `MCPWM5F_IN, `ADCSOC1_IN, `RGMII2RXCTL_IN, 1'b0};
assign input_func_concat_DP6_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS4_IN, `OUTPUTXBAR2_IN, `EPWM1A_IN, `MSC1CLK_IN, `MCPWM4A_IN, `MCPWM8A_IN, `FSI2RXCLK_IN, `MMC0CLK_IN, 1'b0};
assign input_func_concat_DP6_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS5_IN, `OUTPUTXBAR3_IN, `EPWM1B_IN, `MSC1SI_IN, `MCPWM4B_IN, `MCPWM8B_IN, `FSI2RXD0_IN, `MMC0CMD_IN, 1'b0};
assign input_func_concat_DP6_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR4_IN, `EPWM2A_IN, `MSC1SO_IN, `MCPWM4C_IN, `MCPWM8C_IN, `FSI2RXD1_IN, `MMC0DATA0_IN, 1'b0};
assign input_func_concat_DP6_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `OUTPUTXBAR5_IN, `EPWM2B_IN, `MSC1CS0_IN, `MCPWM4D_IN, `MCPWM8D_IN, `FSI3TXCLK_IN, `MMC0DATA1_IN, 1'b0};
assign input_func_concat_DP7_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS4_IN, `SPI2CS4_IN, `MCPWM7E_IN, `MSC0CLK_IN, `LPD_CAN0TX_IN, `LPD_A_PWM1A_IN, 1'b0};
assign input_func_concat_DP7_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI6CS5_IN, `SPI2CS5_IN, `MCPWM7F_IN, `MSC0SI_IN, `LPD_CAN0RX_IN, `LPD_A_PWM1B_IN, 1'b0};
assign input_func_concat_DP7_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM9C_IN, `PSI5_1_RX_IN, `nan_IN, `SDFM8CLK_IN, 1'b0};
assign input_func_concat_DP7_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN9TX_IN, `MCPWM9D_IN, `nan_IN, `SPI8CS4_IN, `SDFM8DATA_IN, 1'b0};
assign input_func_concat_DP7_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN9RX_IN, `MCPWM9E_IN, `nan_IN, `SPI8CS5_IN, `SDFM9CLK_IN, 1'b0};
assign input_func_concat_DP7_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN10TX_IN, `MCPWM9F_IN, `nan_IN, `FSI3RXCLK_IN, `SDFM9DATA_IN, 1'b0};
assign input_func_concat_DP7_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN10RX_IN, `MCPWM10A_IN, `nan_IN, `FSI3RXD0_IN, `SDFM10CLK_IN, 1'b0};
assign input_func_concat_DP7_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MCPWM10B_IN, `nan_IN, `FSI3RXD1_IN, `SDFM10DATA_IN, 1'b0};
assign input_func_concat_DP7_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS4_IN, `EPWM21A_IN, `MCPWM8A_IN, `MSC0SO_IN, `LPD_B_PWM4A_IN, `LPD_A_PWM2A_IN, 1'b0};
assign input_func_concat_DP7_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS5_IN, `EPWM21B_IN, `MCPWM8B_IN, `MSC0CS0_IN, `LPD_B_PWM4B_IN, `LPD_A_PWM2B_IN, 1'b0};
assign input_func_concat_DP7_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS4_IN, `EPWM22A_IN, `MCPWM8C_IN, `MSC0CS1_IN, `LPD_A_PWM1A_IN, `LPD_B_PWM3A_IN, 1'b0};
assign input_func_concat_DP7_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS5_IN, `EPWM22B_IN, `MCPWM8D_IN, `MSC0CS2_IN, `LPD_A_PWM1B_IN, `LPD_B_PWM3B_IN, 1'b0};
assign input_func_concat_DP7_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS4_IN, `EPWM23A_IN, `MCPWM8E_IN, `MSC0CS3_IN, `LPD_A_PWM2A_IN, `LPD_B_PWM4A_IN, 1'b0};
assign input_func_concat_DP7_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI5CS5_IN, `EPWM23B_IN, `MCPWM8F_IN, `PSI5_0_TX_IN, `LPD_A_PWM2B_IN, `LPD_B_PWM4B_IN, 1'b0};
assign input_func_concat_DP7_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM24A_IN, `MCPWM9A_IN, `PSI5_0_RX_IN, `LPD_B_PWM3A_IN, `LPD_CAN0TX_IN, 1'b0};
assign input_func_concat_DP7_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `EPWM24B_IN, `MCPWM9B_IN, `PSI5_1_TX_IN, `LPD_B_PWM3B_IN, `LPD_CAN0RX_IN, 1'b0};
assign input_func_concat_MP0_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS7_IN, `MIBSPI1CS4_IN, `CAN8TX_IN, `SDFM0CLK_IN, 1'b0};
assign input_func_concat_MP0_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS8_IN, `MIBSPI1CS5_IN, `CAN8RX_IN, `SDFM0DATA_IN, 1'b0};
assign input_func_concat_MP0_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS5_IN, `SDFM6CLK_IN, `LIN1TX_IN, `CAN7TX_IN, 1'b0};
assign input_func_concat_MP0_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SDFM6DATA_IN, `LIN1RX_IN, `CAN7RX_IN, 1'b0};
assign input_func_concat_MP0_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS4_IN, `SDFM8CLK_IN, `LIN2TX_IN, `CAN8TX_IN, 1'b0};
assign input_func_concat_MP0_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI4CS5_IN, `SDFM8DATA_IN, `LIN2RX_IN, `CAN8RX_IN, 1'b0};
assign input_func_concat_MP0_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN1TX_IN, `SPI4CS4_IN, `SPI3CS4_IN, `CAN9TX_IN, 1'b0};
assign input_func_concat_MP0_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN1RX_IN, `SPI4CS5_IN, `SPI3CS5_IN, `CAN9RX_IN, 1'b0};
assign input_func_concat_MP0_16 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS5_IN, `nan_IN, `MIBSPI0CS10_IN, `LIN4TX_IN, `CAN10TX_IN, 1'b0};
assign input_func_concat_MP0_17 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN4RX_IN, `CAN10RX_IN, 1'b0};
assign input_func_concat_MP0_18 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS4_IN, `MIBSPI0CS0_IN, `LIN5TX_IN, `CAN11TX_IN, 1'b0};
assign input_func_concat_MP0_19 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS5_IN, `MIBSPI0CS1_IN, `LIN5RX_IN, `CAN11RX_IN, 1'b0};
assign input_func_concat_MP0_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS9_IN, `MIBSPI1CS6_IN, `CAN9TX_IN, `SDFM1CLK_IN, 1'b0};
assign input_func_concat_MP0_20 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN3TX_IN, `MIBSPI0CS2_IN, `LIN6TX_IN, `SPI5CS4_IN, 1'b0};
assign input_func_concat_MP0_21 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN3RX_IN, `MIBSPI0CS3_IN, `LIN6RX_IN, `SPI5CS5_IN, 1'b0};
assign input_func_concat_MP0_22 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS4_IN, `LIN7TX_IN, `SPI6CS4_IN, 1'b0};
assign input_func_concat_MP0_23 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN7RX_IN, `SPI6CS5_IN, 1'b0};
assign input_func_concat_MP0_24 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C0SDA_IN, `SDFM9CLK_IN, `UART0TX_IN, `SDFM11CLK_IN, 1'b0};
assign input_func_concat_MP0_25 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C0SCL_IN, `SDFM9DATA_IN, `UART0RX_IN, `SDFM11DATA_IN, 1'b0};
assign input_func_concat_MP0_26 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C1SDA_IN, `SDFM10CLK_IN, `UART1TX_IN, `LIN4TX_IN, 1'b0};
assign input_func_concat_MP0_27 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C1SCL_IN, `SDFM10DATA_IN, `UART1RX_IN, `LIN4RX_IN, 1'b0};
assign input_func_concat_MP0_28 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS11_IN, `LIN3TX_IN, `LIN5TX_IN, 1'b0};
assign input_func_concat_MP0_29 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `LIN3RX_IN, `LIN5RX_IN, 1'b0};
assign input_func_concat_MP0_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS10_IN, `MIBSPI1CS7_IN, `CAN9RX_IN, `SDFM1DATA_IN, 1'b0};
assign input_func_concat_MP0_30 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C2SDA_IN, `MIBSPI0CS5_IN, `SPI6CS4_IN, `LIN6TX_IN, 1'b0};
assign input_func_concat_MP0_31 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C2SCL_IN, `MIBSPI0CS6_IN, `SPI6CS5_IN, `LIN6RX_IN, 1'b0};
assign input_func_concat_MP0_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS11_IN, `MIBSPI1CS8_IN, `CAN10TX_IN, `SDFM2CLK_IN, 1'b0};
assign input_func_concat_MP0_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN10RX_IN, `SDFM2DATA_IN, 1'b0};
assign input_func_concat_MP0_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI8CS4_IN, `MIBSPI1CS9_IN, `CAN11TX_IN, `SDFM3CLK_IN, 1'b0};
assign input_func_concat_MP0_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI8CS5_IN, `MIBSPI1CS10_IN, `CAN11RX_IN, `SDFM3DATA_IN, 1'b0};
assign input_func_concat_MP0_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI9CS4_IN, `MIBSPI1CS11_IN, `SDFM5CLK_IN, `LIN0TX_IN, `CAN6TX_IN, 1'b0};
assign input_func_concat_MP0_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS4_IN, `SDFM5DATA_IN, `LIN0RX_IN, `CAN6RX_IN, 1'b0};
assign input_func_concat_MP1_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C3SDA_IN, `MIBSPI0CS7_IN, `SPI7CS4_IN, `LIN7TX_IN, 1'b0};
assign input_func_concat_MP1_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `I2C3SCL_IN, `MIBSPI0CS8_IN, `SPI7CS5_IN, `LIN7RX_IN, 1'b0};
assign input_func_concat_MP1_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS10_IN, `SPI5CS4_IN, 1'b0};
assign input_func_concat_MP1_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS11_IN, `SPI5CS5_IN, 1'b0};
assign input_func_concat_MP1_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS4_IN, 1'b0};
assign input_func_concat_MP1_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS5_IN, 1'b0};
assign input_func_concat_MP1_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS6_IN, 1'b0};
assign input_func_concat_MP1_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS7_IN, 1'b0};
assign input_func_concat_MP1_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI0CS9_IN, `SENT4TXRX_IN, `UART1TX_IN, 1'b0};
assign input_func_concat_MP1_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SENT5TXRX_IN, `UART1RX_IN, 1'b0};
assign input_func_concat_MP1_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS4_IN, `SENT0TXRX_IN, 1'b0};
assign input_func_concat_MP1_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS5_IN, `SENT1TXRX_IN, 1'b0};
assign input_func_concat_MP1_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS6_IN, `SENT2TXRX_IN, 1'b0};
assign input_func_concat_MP1_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS7_IN, `SENT3TXRX_IN, 1'b0};
assign input_func_concat_MP1_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS8_IN, `SENT4TXRX_IN, 1'b0};
assign input_func_concat_MP1_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS9_IN, `SENT5TXRX_IN, 1'b0};
assign input_func_concat_MP2_0 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN11TX_IN, `MCPWM10C_IN, `I2C0SDA_IN, `CAN0TX_IN, `SDFM4CLK_IN, 1'b0};
assign input_func_concat_MP2_1 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `CAN11RX_IN, `MCPWM10D_IN, `I2C0SCL_IN, `CAN0RX_IN, `SDFM4DATA_IN, 1'b0};
assign input_func_concat_MP2_10 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS1_IN, `SDFM2CLK_IN, `CAN5TX_IN, `SPI6CS4_IN, 1'b0};
assign input_func_concat_MP2_11 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS2_IN, `SDFM2DATA_IN, `CAN5RX_IN, `SPI6CS5_IN, 1'b0};
assign input_func_concat_MP2_12 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS3_IN, `SDFM3CLK_IN, `CAN6TX_IN, `SENT4TXRX_IN, 1'b0};
assign input_func_concat_MP2_13 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS4_IN, `SDFM3DATA_IN, `CAN6RX_IN, `SENT5TXRX_IN, 1'b0};
assign input_func_concat_MP2_14 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS5_IN, `SDFM4CLK_IN, `CAN7TX_IN, `LPD_LIN0TX_IN, 1'b0};
assign input_func_concat_MP2_15 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS6_IN, `SDFM4DATA_IN, `CAN7RX_IN, `LPD_LIN0RX_IN, 1'b0};
assign input_func_concat_MP2_2 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS4_IN, `MCPWM10E_IN, `I2C1SDA_IN, `CAN1TX_IN, `SDFM5CLK_IN, 1'b0};
assign input_func_concat_MP2_3 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SPI7CS5_IN, `MCPWM10F_IN, `I2C1SCL_IN, `CAN1RX_IN, `SDFM5DATA_IN, 1'b0};
assign input_func_concat_MP2_4 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `RDC0PWM_N_IN, `SPI3CS4_IN, `I2C2SDA_IN, `CAN2TX_IN, `SDFM6CLK_IN, 1'b0};
assign input_func_concat_MP2_5 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `RDC0PWM_P_IN, `SPI3CS5_IN, `I2C2SCL_IN, `CAN2RX_IN, `SDFM6DATA_IN, 1'b0};
assign input_func_concat_MP2_6 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `RDC1PWM_N_IN, `SPI8CS4_IN, `I2C3SDA_IN, `CAN3TX_IN, `SDFM7CLK_IN, 1'b0};
assign input_func_concat_MP2_7 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `RDC1PWM_P_IN, `SPI8CS5_IN, `I2C3SCL_IN, `CAN3RX_IN, `SDFM7DATA_IN, 1'b0};
assign input_func_concat_MP2_8 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `SDFM1CLK_IN, `CAN4TX_IN, `LPD_LIN0TX_IN, 1'b0};
assign input_func_concat_MP2_9 = {`nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `nan_IN, `MIBSPI1CS0_IN, `SDFM1DATA_IN, `CAN4RX_IN, `LPD_LIN0RX_IN, 1'b0};
assign nan_IN = 1'b0;

// Properties
 property iomux_output_drive(logic funcsel, logic gpioouten, logic oe, logic od, logic func_out, logic pad);
  (funcsel == 1 && gpioouten == 1 && oe == 1 && od == 0) |-> (pad == func_out);
 endproperty
 property iomux_output_open_drain(logic funcsel, logic gpioouten, logic oe, logic od, logic func_out, logic pad, logic pad_gz);
  (funcsel == 1 && gpioouten == 1 && oe == 1 && od == 1) |-> (pad_gz == !func_out && pad == 0);
 endproperty
 property iomux_pull_up(logic pullen, logic pullsel, logic pad_pullup);
  (pullen == 1 && pullsel == `PULL_UP) |-> (pad_pullup == 1);
 endproperty
 property iomux_pull_up_reverse(logic pad_pullup, logic pullen, logic pullsel);
  (pad_pullup == 1) |-> (pullen == 1 && pullsel == `PULL_UP);
 endproperty
 property iomux_pull_down(logic pullen, logic pullsel, logic pad_pd);
  (pullen == 1 && pullsel == `PULL_DOWN) |-> (pad_pd == 0);
 endproperty
 property iomux_pull_down_reverse(logic pad_pd, logic pullen, logic pullsel);
  (pad_pd == 0) |-> (pullen == 1 && pullsel == `PULL_DOWN);
 endproperty
 property iomux_highz_conditions(logic pullen, logic outen, logic pad);
  (pullen == 0 && outen == 0) |-> (pad == 1'bz);
 endproperty
 property iomux_highz_reverse(logic pad, logic pullen, logic outen);
  (pad == 1'bz) |-> (pullen == 0 && outen == 0);
 endproperty
 property iomux_input_path(logic ie, logic outen, logic [31:0] infunc_en, logic [31:0] in_concat, logic [31:0] pad, logic [31:0] default_value);
  (ie == 1 && outen == 0) |-> (in_concat == (infunc_en & {32{pad}}) | ~infunc_en & {default_value});
 endproperty

// Assertions
ap_DP0_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_0),
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE)
));
ap_DP0_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_0_PINCTRL_0_IE),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_0),
  .pad(`DP0_0),
  .default_value(`default_value)));
ap_DP0_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCLK_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`TPIUCLK_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCLK_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`TPIUCLK_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_0),
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE)
));
ap_DP0_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_0_PINCTRL_0_IE),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_0),
  .pad(`DP0_0),
  .default_value(`default_value)));
ap_DP0_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_0_OUTFUNC_SEL),
  .gpioouten(`DP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP0_0_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP0_0),
  .pad_gz(`DP0_0_pad_y)
));
ap_DP0_0_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_0)
));
ap_DP0_0_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_0),
  .pullen(`DP0_0_PULLEN),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE)
));
ap_DP0_0_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_0_PINCTRL_0_IE),
  .outen(`DP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_0),
  .pad(`DP0_0),
  .default_value(`default_value)));
ap_DP0_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_0_PULLEN),
  .pullsel(`DP0_0_PULLSEL),
  .pad_pullup(`DP0_0)
));
ap_DP0_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_0),
  .pullen(`DP0_0_PULLEN),
  .pullsel(`DP0_0_PULLSEL)
));
ap_DP0_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_0_PULLEN),
  .pullsel(`DP0_0_PULLSEL),
  .pad_pd(`DP0_0)
));
ap_DP0_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_0),
  .pullen(`DP0_0_PULLEN),
  .pullsel(`DP0_0_PULLSEL)
));
ap_DP0_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_1),
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE)
));
ap_DP0_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_1_PINCTRL_0_IE),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_1),
  .pad(`DP0_1),
  .default_value(`default_value)));
ap_DP0_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCTL_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`TPIUCTL_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCTL_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`TPIUCTL_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_1),
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE)
));
ap_DP0_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_1_PINCTRL_0_IE),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_1),
  .pad(`DP0_1),
  .default_value(`default_value)));
ap_DP0_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_1_OUTFUNC_SEL),
  .gpioouten(`DP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP0_1_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP0_1),
  .pad_gz(`DP0_1_pad_y)
));
ap_DP0_1_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_1)
));
ap_DP0_1_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_1),
  .pullen(`DP0_1_PULLEN),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE)
));
ap_DP0_1_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_1_PINCTRL_0_IE),
  .outen(`DP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_1),
  .pad(`DP0_1),
  .default_value(`default_value)));
ap_DP0_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_1_PULLEN),
  .pullsel(`DP0_1_PULLSEL),
  .pad_pullup(`DP0_1)
));
ap_DP0_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_1),
  .pullen(`DP0_1_PULLEN),
  .pullsel(`DP0_1_PULLSEL)
));
ap_DP0_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_1_PULLEN),
  .pullsel(`DP0_1_PULLSEL),
  .pad_pd(`DP0_1)
));
ap_DP0_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_1),
  .pullen(`DP0_1_PULLEN),
  .pullsel(`DP0_1_PULLSEL)
));
ap_DP0_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_2),
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE)
));
ap_DP0_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_2_PINCTRL_0_IE),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_2),
  .pad(`DP0_2),
  .default_value(`default_value)));
ap_DP0_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA0_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`TPIUDATA0_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA0_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`TPIUDATA0_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_2),
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE)
));
ap_DP0_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_2_PINCTRL_0_IE),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_2),
  .pad(`DP0_2),
  .default_value(`default_value)));
ap_DP0_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_2_OUTFUNC_SEL),
  .gpioouten(`DP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP0_2_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP0_2),
  .pad_gz(`DP0_2_pad_y)
));
ap_DP0_2_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_2)
));
ap_DP0_2_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_2),
  .pullen(`DP0_2_PULLEN),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE)
));
ap_DP0_2_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_2_PINCTRL_0_IE),
  .outen(`DP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_2),
  .pad(`DP0_2),
  .default_value(`default_value)));
ap_DP0_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_2_PULLEN),
  .pullsel(`DP0_2_PULLSEL),
  .pad_pullup(`DP0_2)
));
ap_DP0_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_2),
  .pullen(`DP0_2_PULLEN),
  .pullsel(`DP0_2_PULLSEL)
));
ap_DP0_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_2_PULLEN),
  .pullsel(`DP0_2_PULLSEL),
  .pad_pd(`DP0_2)
));
ap_DP0_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_2),
  .pullen(`DP0_2_PULLEN),
  .pullsel(`DP0_2_PULLSEL)
));
ap_DP0_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_3),
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE)
));
ap_DP0_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_3_PINCTRL_0_IE),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_3),
  .pad(`DP0_3),
  .default_value(`default_value)));
ap_DP0_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA1_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`TPIUDATA1_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA1_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`TPIUDATA1_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_3),
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE)
));
ap_DP0_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_3_PINCTRL_0_IE),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_3),
  .pad(`DP0_3),
  .default_value(`default_value)));
ap_DP0_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_3_OUTFUNC_SEL),
  .gpioouten(`DP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP0_3_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP0_3),
  .pad_gz(`DP0_3_pad_y)
));
ap_DP0_3_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_3)
));
ap_DP0_3_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_3),
  .pullen(`DP0_3_PULLEN),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE)
));
ap_DP0_3_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_3_PINCTRL_0_IE),
  .outen(`DP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_3),
  .pad(`DP0_3),
  .default_value(`default_value)));
ap_DP0_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_3_PULLEN),
  .pullsel(`DP0_3_PULLSEL),
  .pad_pullup(`DP0_3)
));
ap_DP0_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_3),
  .pullen(`DP0_3_PULLEN),
  .pullsel(`DP0_3_PULLSEL)
));
ap_DP0_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_3_PULLEN),
  .pullsel(`DP0_3_PULLSEL),
  .pad_pd(`DP0_3)
));
ap_DP0_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_3),
  .pullen(`DP0_3_PULLEN),
  .pullsel(`DP0_3_PULLSEL)
));
ap_DP0_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_4),
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE)
));
ap_DP0_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_4_PINCTRL_0_IE),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_4),
  .pad(`DP0_4),
  .default_value(`default_value)));
ap_DP0_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA2_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`TPIUDATA2_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA2_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`TPIUDATA2_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_4),
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE)
));
ap_DP0_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_4_PINCTRL_0_IE),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_4),
  .pad(`DP0_4),
  .default_value(`default_value)));
ap_DP0_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_4_OUTFUNC_SEL),
  .gpioouten(`DP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP0_4_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP0_4),
  .pad_gz(`DP0_4_pad_y)
));
ap_DP0_4_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_4)
));
ap_DP0_4_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_4),
  .pullen(`DP0_4_PULLEN),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE)
));
ap_DP0_4_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_4_PINCTRL_0_IE),
  .outen(`DP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_4),
  .pad(`DP0_4),
  .default_value(`default_value)));
ap_DP0_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_4_PULLEN),
  .pullsel(`DP0_4_PULLSEL),
  .pad_pullup(`DP0_4)
));
ap_DP0_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_4),
  .pullen(`DP0_4_PULLEN),
  .pullsel(`DP0_4_PULLSEL)
));
ap_DP0_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_4_PULLEN),
  .pullsel(`DP0_4_PULLSEL),
  .pad_pd(`DP0_4)
));
ap_DP0_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_4),
  .pullen(`DP0_4_PULLEN),
  .pullsel(`DP0_4_PULLSEL)
));
ap_DP0_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_5),
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE)
));
ap_DP0_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_5_PINCTRL_0_IE),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_5),
  .pad(`DP0_5),
  .default_value(`default_value)));
ap_DP0_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA3_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`TPIUDATA3_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA3_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`TPIUDATA3_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_5),
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE)
));
ap_DP0_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_5_PINCTRL_0_IE),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_5),
  .pad(`DP0_5),
  .default_value(`default_value)));
ap_DP0_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_5_OUTFUNC_SEL),
  .gpioouten(`DP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP0_5_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP0_5),
  .pad_gz(`DP0_5_pad_y)
));
ap_DP0_5_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_5)
));
ap_DP0_5_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_5),
  .pullen(`DP0_5_PULLEN),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE)
));
ap_DP0_5_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_5_PINCTRL_0_IE),
  .outen(`DP0_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_5),
  .pad(`DP0_5),
  .default_value(`default_value)));
ap_DP0_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_5_PULLEN),
  .pullsel(`DP0_5_PULLSEL),
  .pad_pullup(`DP0_5)
));
ap_DP0_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_5),
  .pullen(`DP0_5_PULLEN),
  .pullsel(`DP0_5_PULLSEL)
));
ap_DP0_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_5_PULLEN),
  .pullsel(`DP0_5_PULLSEL),
  .pad_pd(`DP0_5)
));
ap_DP0_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_5),
  .pullen(`DP0_5_PULLEN),
  .pullsel(`DP0_5_PULLSEL)
));
ap_DP0_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_6),
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE)
));
ap_DP0_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_6_PINCTRL_0_IE),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_6),
  .pad(`DP0_6),
  .default_value(`default_value)));
ap_DP0_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_6),
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE)
));
ap_DP0_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_6_PINCTRL_0_IE),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_6),
  .pad(`DP0_6),
  .default_value(`default_value)));
ap_DP0_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_6_OUTFUNC_SEL),
  .gpioouten(`DP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP0_6_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP0_6),
  .pad_gz(`DP0_6_pad_y)
));
ap_DP0_6_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_6)
));
ap_DP0_6_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_6),
  .pullen(`DP0_6_PULLEN),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE)
));
ap_DP0_6_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_6_PINCTRL_0_IE),
  .outen(`DP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_6),
  .pad(`DP0_6),
  .default_value(`default_value)));
ap_DP0_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_6_PULLEN),
  .pullsel(`DP0_6_PULLSEL),
  .pad_pullup(`DP0_6)
));
ap_DP0_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_6),
  .pullen(`DP0_6_PULLEN),
  .pullsel(`DP0_6_PULLSEL)
));
ap_DP0_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_6_PULLEN),
  .pullsel(`DP0_6_PULLSEL),
  .pad_pd(`DP0_6)
));
ap_DP0_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_6),
  .pullen(`DP0_6_PULLEN),
  .pullsel(`DP0_6_PULLSEL)
));
ap_DP0_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_7),
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE)
));
ap_DP0_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_7_PINCTRL_0_IE),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_7),
  .pad(`DP0_7),
  .default_value(`default_value)));
ap_DP0_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_7),
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE)
));
ap_DP0_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_7_PINCTRL_0_IE),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_7),
  .pad(`DP0_7),
  .default_value(`default_value)));
ap_DP0_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_7_OUTFUNC_SEL),
  .gpioouten(`DP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP0_7_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP0_7),
  .pad_gz(`DP0_7_pad_y)
));
ap_DP0_7_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_7)
));
ap_DP0_7_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_7),
  .pullen(`DP0_7_PULLEN),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE)
));
ap_DP0_7_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_7_PINCTRL_0_IE),
  .outen(`DP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_7),
  .pad(`DP0_7),
  .default_value(`default_value)));
ap_DP0_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_7_PULLEN),
  .pullsel(`DP0_7_PULLSEL),
  .pad_pullup(`DP0_7)
));
ap_DP0_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_7),
  .pullen(`DP0_7_PULLEN),
  .pullsel(`DP0_7_PULLSEL)
));
ap_DP0_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_7_PULLEN),
  .pullsel(`DP0_7_PULLSEL),
  .pad_pd(`DP0_7)
));
ap_DP0_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_7),
  .pullen(`DP0_7_PULLEN),
  .pullsel(`DP0_7_PULLSEL)
));
ap_DP0_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_8),
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE)
));
ap_DP0_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_8_PINCTRL_0_IE),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_8),
  .pad(`DP0_8),
  .default_value(`default_value)));
ap_DP0_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_8),
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE)
));
ap_DP0_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_8_PINCTRL_0_IE),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_8),
  .pad(`DP0_8),
  .default_value(`default_value)));
ap_DP0_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_8_OUTFUNC_SEL),
  .gpioouten(`DP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP0_8_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP0_8),
  .pad_gz(`DP0_8_pad_y)
));
ap_DP0_8_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_8)
));
ap_DP0_8_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_8),
  .pullen(`DP0_8_PULLEN),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE)
));
ap_DP0_8_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_8_PINCTRL_0_IE),
  .outen(`DP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_8),
  .pad(`DP0_8),
  .default_value(`default_value)));
ap_DP0_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_8_PULLEN),
  .pullsel(`DP0_8_PULLSEL),
  .pad_pullup(`DP0_8)
));
ap_DP0_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_8),
  .pullen(`DP0_8_PULLEN),
  .pullsel(`DP0_8_PULLSEL)
));
ap_DP0_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_8_PULLEN),
  .pullsel(`DP0_8_PULLSEL),
  .pad_pd(`DP0_8)
));
ap_DP0_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_8),
  .pullen(`DP0_8_PULLEN),
  .pullsel(`DP0_8_PULLSEL)
));
ap_DP0_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_9),
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE)
));
ap_DP0_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_9_PINCTRL_0_IE),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_9),
  .pad(`DP0_9),
  .default_value(`default_value)));
ap_DP0_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_9),
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE)
));
ap_DP0_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_9_PINCTRL_0_IE),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_9),
  .pad(`DP0_9),
  .default_value(`default_value)));
ap_DP0_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_9_OUTFUNC_SEL),
  .gpioouten(`DP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP0_9_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP0_9),
  .pad_gz(`DP0_9_pad_y)
));
ap_DP0_9_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_9)
));
ap_DP0_9_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_9),
  .pullen(`DP0_9_PULLEN),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE)
));
ap_DP0_9_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_9_PINCTRL_0_IE),
  .outen(`DP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_9),
  .pad(`DP0_9),
  .default_value(`default_value)));
ap_DP0_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_9_PULLEN),
  .pullsel(`DP0_9_PULLSEL),
  .pad_pullup(`DP0_9)
));
ap_DP0_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_9),
  .pullen(`DP0_9_PULLEN),
  .pullsel(`DP0_9_PULLSEL)
));
ap_DP0_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_9_PULLEN),
  .pullsel(`DP0_9_PULLSEL),
  .pad_pd(`DP0_9)
));
ap_DP0_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_9),
  .pullen(`DP0_9_PULLEN),
  .pullsel(`DP0_9_PULLSEL)
));
ap_DP0_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXCLK_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`FSI0TXCLK_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXCLK_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`FSI0TXCLK_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE)
));
ap_DP0_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_10_PINCTRL_0_IE),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_10),
  .pad(`DP0_10),
  .default_value(`default_value)));
ap_DP0_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE)
));
ap_DP0_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_10_PINCTRL_0_IE),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_10),
  .pad(`DP0_10),
  .default_value(`default_value)));
ap_DP0_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE)
));
ap_DP0_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_10_PINCTRL_0_IE),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_10),
  .pad(`DP0_10),
  .default_value(`default_value)));
ap_DP0_10_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_10_OUTFUNC_SEL),
  .gpioouten(`DP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP0_10_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP0_10),
  .pad_gz(`DP0_10_pad_y)
));
ap_DP0_10_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_10)
));
ap_DP0_10_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE)
));
ap_DP0_10_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_10_PINCTRL_0_IE),
  .outen(`DP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_10),
  .pad(`DP0_10),
  .default_value(`default_value)));
ap_DP0_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_10_PULLEN),
  .pullsel(`DP0_10_PULLSEL),
  .pad_pullup(`DP0_10)
));
ap_DP0_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .pullsel(`DP0_10_PULLSEL)
));
ap_DP0_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_10_PULLEN),
  .pullsel(`DP0_10_PULLSEL),
  .pad_pd(`DP0_10)
));
ap_DP0_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_10),
  .pullen(`DP0_10_PULLEN),
  .pullsel(`DP0_10_PULLSEL)
));
ap_DP0_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD0_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`FSI0TXD0_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD0_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`FSI0TXD0_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE)
));
ap_DP0_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_11_PINCTRL_0_IE),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_11),
  .pad(`DP0_11),
  .default_value(`default_value)));
ap_DP0_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE)
));
ap_DP0_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_11_PINCTRL_0_IE),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_11),
  .pad(`DP0_11),
  .default_value(`default_value)));
ap_DP0_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE)
));
ap_DP0_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_11_PINCTRL_0_IE),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_11),
  .pad(`DP0_11),
  .default_value(`default_value)));
ap_DP0_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_11_OUTFUNC_SEL),
  .gpioouten(`DP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP0_11_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP0_11),
  .pad_gz(`DP0_11_pad_y)
));
ap_DP0_11_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_11)
));
ap_DP0_11_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE)
));
ap_DP0_11_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_11_PINCTRL_0_IE),
  .outen(`DP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_11),
  .pad(`DP0_11),
  .default_value(`default_value)));
ap_DP0_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_11_PULLEN),
  .pullsel(`DP0_11_PULLSEL),
  .pad_pullup(`DP0_11)
));
ap_DP0_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .pullsel(`DP0_11_PULLSEL)
));
ap_DP0_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_11_PULLEN),
  .pullsel(`DP0_11_PULLSEL),
  .pad_pd(`DP0_11)
));
ap_DP0_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_11),
  .pullen(`DP0_11_PULLEN),
  .pullsel(`DP0_11_PULLSEL)
));
ap_DP0_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD1_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`FSI0TXD1_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD1_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`FSI0TXD1_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE)
));
ap_DP0_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_12_PINCTRL_0_IE),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_12),
  .pad(`DP0_12),
  .default_value(`default_value)));
ap_DP0_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE)
));
ap_DP0_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_12_PINCTRL_0_IE),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_12),
  .pad(`DP0_12),
  .default_value(`default_value)));
ap_DP0_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE)
));
ap_DP0_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_12_PINCTRL_0_IE),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_12),
  .pad(`DP0_12),
  .default_value(`default_value)));
ap_DP0_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_12_OUTFUNC_SEL),
  .gpioouten(`DP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP0_12_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP0_12),
  .pad_gz(`DP0_12_pad_y)
));
ap_DP0_12_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_12)
));
ap_DP0_12_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE)
));
ap_DP0_12_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_12_PINCTRL_0_IE),
  .outen(`DP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_12),
  .pad(`DP0_12),
  .default_value(`default_value)));
ap_DP0_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_12_PULLEN),
  .pullsel(`DP0_12_PULLSEL),
  .pad_pullup(`DP0_12)
));
ap_DP0_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .pullsel(`DP0_12_PULLSEL)
));
ap_DP0_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_12_PULLEN),
  .pullsel(`DP0_12_PULLSEL),
  .pad_pd(`DP0_12)
));
ap_DP0_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_12),
  .pullen(`DP0_12_PULLEN),
  .pullsel(`DP0_12_PULLSEL)
));
ap_DP0_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXCLK_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`FSI0RXCLK_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXCLK_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`FSI0RXCLK_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE)
));
ap_DP0_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_13_PINCTRL_0_IE),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_13),
  .pad(`DP0_13),
  .default_value(`default_value)));
ap_DP0_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE)
));
ap_DP0_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_13_PINCTRL_0_IE),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_13),
  .pad(`DP0_13),
  .default_value(`default_value)));
ap_DP0_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXCLK_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`FSI0TXCLK_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXCLK_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`FSI0TXCLK_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE)
));
ap_DP0_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_13_PINCTRL_0_IE),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_13),
  .pad(`DP0_13),
  .default_value(`default_value)));
ap_DP0_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE)
));
ap_DP0_13_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_13_PINCTRL_0_IE),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_13),
  .pad(`DP0_13),
  .default_value(`default_value)));
ap_DP0_13_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_13_OUTFUNC_SEL),
  .gpioouten(`DP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP0_13_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP0_13),
  .pad_gz(`DP0_13_pad_y)
));
ap_DP0_13_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_13)
));
ap_DP0_13_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE)
));
ap_DP0_13_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_13_PINCTRL_0_IE),
  .outen(`DP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_13),
  .pad(`DP0_13),
  .default_value(`default_value)));
ap_DP0_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_13_PULLEN),
  .pullsel(`DP0_13_PULLSEL),
  .pad_pullup(`DP0_13)
));
ap_DP0_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .pullsel(`DP0_13_PULLSEL)
));
ap_DP0_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_13_PULLEN),
  .pullsel(`DP0_13_PULLSEL),
  .pad_pd(`DP0_13)
));
ap_DP0_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_13),
  .pullen(`DP0_13_PULLEN),
  .pullsel(`DP0_13_PULLSEL)
));
ap_DP0_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD0_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`FSI0RXD0_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD0_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`FSI0RXD0_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD0_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`FSI0TXD0_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD0_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`FSI0TXD0_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_14_OUTFUNC_SEL),
  .gpioouten(`DP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP0_14_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP0_14),
  .pad_gz(`DP0_14_pad_y)
));
ap_DP0_14_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_14)
));
ap_DP0_14_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE)
));
ap_DP0_14_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_14_PINCTRL_0_IE),
  .outen(`DP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_14),
  .pad(`DP0_14),
  .default_value(`default_value)));
ap_DP0_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_14_PULLEN),
  .pullsel(`DP0_14_PULLSEL),
  .pad_pullup(`DP0_14)
));
ap_DP0_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .pullsel(`DP0_14_PULLSEL)
));
ap_DP0_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_14_PULLEN),
  .pullsel(`DP0_14_PULLSEL),
  .pad_pd(`DP0_14)
));
ap_DP0_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_14),
  .pullen(`DP0_14_PULLEN),
  .pullsel(`DP0_14_PULLSEL)
));
ap_DP0_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD1_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`FSI0RXD1_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD1_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`FSI0RXD1_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD1_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`FSI0TXD1_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0TXD1_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`FSI0TXD1_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_15_OUTFUNC_SEL),
  .gpioouten(`DP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP0_15_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP0_15),
  .pad_gz(`DP0_15_pad_y)
));
ap_DP0_15_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_15)
));
ap_DP0_15_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE)
));
ap_DP0_15_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_15_PINCTRL_0_IE),
  .outen(`DP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_15),
  .pad(`DP0_15),
  .default_value(`default_value)));
ap_DP0_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_15_PULLEN),
  .pullsel(`DP0_15_PULLSEL),
  .pad_pullup(`DP0_15)
));
ap_DP0_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .pullsel(`DP0_15_PULLSEL)
));
ap_DP0_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_15_PULLEN),
  .pullsel(`DP0_15_PULLSEL),
  .pad_pd(`DP0_15)
));
ap_DP0_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_15),
  .pullen(`DP0_15_PULLEN),
  .pullsel(`DP0_15_PULLSEL)
));
ap_DP0_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE)
));
ap_DP0_16_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_16_PINCTRL_0_IE),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_16),
  .pad(`DP0_16),
  .default_value(`default_value)));
ap_DP0_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXCLK_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`FSI0RXCLK_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXCLK_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`FSI0RXCLK_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE)
));
ap_DP0_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_16_PINCTRL_0_IE),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_16),
  .pad(`DP0_16),
  .default_value(`default_value)));
ap_DP0_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE)
));
ap_DP0_16_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_16_PINCTRL_0_IE),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_16),
  .pad(`DP0_16),
  .default_value(`default_value)));
ap_DP0_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE)
));
ap_DP0_16_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_16_PINCTRL_0_IE),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_16),
  .pad(`DP0_16),
  .default_value(`default_value)));
ap_DP0_16_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_16_OUTFUNC_SEL),
  .gpioouten(`DP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP0_16_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP0_16),
  .pad_gz(`DP0_16_pad_y)
));
ap_DP0_16_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_16)
));
ap_DP0_16_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE)
));
ap_DP0_16_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_16_PINCTRL_0_IE),
  .outen(`DP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_16),
  .pad(`DP0_16),
  .default_value(`default_value)));
ap_DP0_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_16_PULLEN),
  .pullsel(`DP0_16_PULLSEL),
  .pad_pullup(`DP0_16)
));
ap_DP0_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .pullsel(`DP0_16_PULLSEL)
));
ap_DP0_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_16_PULLEN),
  .pullsel(`DP0_16_PULLSEL),
  .pad_pd(`DP0_16)
));
ap_DP0_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_16),
  .pullen(`DP0_16_PULLEN),
  .pullsel(`DP0_16_PULLSEL)
));
ap_DP0_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE)
));
ap_DP0_17_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_17_PINCTRL_0_IE),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_17),
  .pad(`DP0_17),
  .default_value(`default_value)));
ap_DP0_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD0_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`FSI0RXD0_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD0_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`FSI0RXD0_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE)
));
ap_DP0_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_17_PINCTRL_0_IE),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_17),
  .pad(`DP0_17),
  .default_value(`default_value)));
ap_DP0_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE)
));
ap_DP0_17_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_17_PINCTRL_0_IE),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_17),
  .pad(`DP0_17),
  .default_value(`default_value)));
ap_DP0_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE)
));
ap_DP0_17_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_17_PINCTRL_0_IE),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_17),
  .pad(`DP0_17),
  .default_value(`default_value)));
ap_DP0_17_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_17_OUTFUNC_SEL),
  .gpioouten(`DP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP0_17_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP0_17),
  .pad_gz(`DP0_17_pad_y)
));
ap_DP0_17_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_17)
));
ap_DP0_17_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE)
));
ap_DP0_17_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_17_PINCTRL_0_IE),
  .outen(`DP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_17),
  .pad(`DP0_17),
  .default_value(`default_value)));
ap_DP0_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_17_PULLEN),
  .pullsel(`DP0_17_PULLSEL),
  .pad_pullup(`DP0_17)
));
ap_DP0_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .pullsel(`DP0_17_PULLSEL)
));
ap_DP0_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_17_PULLEN),
  .pullsel(`DP0_17_PULLSEL),
  .pad_pd(`DP0_17)
));
ap_DP0_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_17),
  .pullen(`DP0_17_PULLEN),
  .pullsel(`DP0_17_PULLSEL)
));
ap_DP0_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD1_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`FSI0RXD1_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`FSI0RXD1_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`FSI0RXD1_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_18_OUTFUNC_SEL),
  .gpioouten(`DP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP0_18_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP0_18),
  .pad_gz(`DP0_18_pad_y)
));
ap_DP0_18_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_18)
));
ap_DP0_18_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE)
));
ap_DP0_18_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_18_PINCTRL_0_IE),
  .outen(`DP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_18),
  .pad(`DP0_18),
  .default_value(`default_value)));
ap_DP0_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_18_PULLEN),
  .pullsel(`DP0_18_PULLSEL),
  .pad_pullup(`DP0_18)
));
ap_DP0_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .pullsel(`DP0_18_PULLSEL)
));
ap_DP0_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_18_PULLEN),
  .pullsel(`DP0_18_PULLSEL),
  .pad_pd(`DP0_18)
));
ap_DP0_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_18),
  .pullen(`DP0_18_PULLEN),
  .pullsel(`DP0_18_PULLSEL)
));
ap_DP0_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_19_OUTFUNC_SEL),
  .gpioouten(`DP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP0_19_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP0_19),
  .pad_gz(`DP0_19_pad_y)
));
ap_DP0_19_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_19)
));
ap_DP0_19_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE)
));
ap_DP0_19_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP0_19_PINCTRL_0_IE),
  .outen(`DP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_19),
  .pad(`DP0_19),
  .default_value(`default_value)));
ap_DP0_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_19_PULLEN),
  .pullsel(`DP0_19_PULLSEL),
  .pad_pullup(`DP0_19)
));
ap_DP0_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .pullsel(`DP0_19_PULLSEL)
));
ap_DP0_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_19_PULLEN),
  .pullsel(`DP0_19_PULLSEL),
  .pad_pd(`DP0_19)
));
ap_DP0_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_19),
  .pullen(`DP0_19_PULLEN),
  .pullsel(`DP0_19_PULLSEL)
));
ap_DP0_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE)
));
ap_DP0_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_20_PINCTRL_0_IE),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_20),
  .pad(`DP0_20),
  .default_value(`default_value)));
ap_DP0_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE)
));
ap_DP0_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_20_PINCTRL_0_IE),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_20),
  .pad(`DP0_20),
  .default_value(`default_value)));
ap_DP0_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE)
));
ap_DP0_20_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_20_PINCTRL_0_IE),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_20),
  .pad(`DP0_20),
  .default_value(`default_value)));
ap_DP0_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_20_OUTFUNC_SEL),
  .gpioouten(`DP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP0_20_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP0_20),
  .pad_gz(`DP0_20_pad_y)
));
ap_DP0_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_20)
));
ap_DP0_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE)
));
ap_DP0_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_20_PINCTRL_0_IE),
  .outen(`DP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_20),
  .pad(`DP0_20),
  .default_value(`default_value)));
ap_DP0_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_20_PULLEN),
  .pullsel(`DP0_20_PULLSEL),
  .pad_pullup(`DP0_20)
));
ap_DP0_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .pullsel(`DP0_20_PULLSEL)
));
ap_DP0_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_20_PULLEN),
  .pullsel(`DP0_20_PULLSEL),
  .pad_pd(`DP0_20)
));
ap_DP0_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_20),
  .pullen(`DP0_20_PULLEN),
  .pullsel(`DP0_20_PULLSEL)
));
ap_DP0_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE)
));
ap_DP0_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_21_PINCTRL_0_IE),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_21),
  .pad(`DP0_21),
  .default_value(`default_value)));
ap_DP0_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE)
));
ap_DP0_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_21_PINCTRL_0_IE),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_21),
  .pad(`DP0_21),
  .default_value(`default_value)));
ap_DP0_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE)
));
ap_DP0_21_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_21_PINCTRL_0_IE),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_21),
  .pad(`DP0_21),
  .default_value(`default_value)));
ap_DP0_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_21_OUTFUNC_SEL),
  .gpioouten(`DP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`DP0_21_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`DP0_21),
  .pad_gz(`DP0_21_pad_y)
));
ap_DP0_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_21)
));
ap_DP0_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE)
));
ap_DP0_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_21_PINCTRL_0_IE),
  .outen(`DP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_21),
  .pad(`DP0_21),
  .default_value(`default_value)));
ap_DP0_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_21_PULLEN),
  .pullsel(`DP0_21_PULLSEL),
  .pad_pullup(`DP0_21)
));
ap_DP0_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .pullsel(`DP0_21_PULLSEL)
));
ap_DP0_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_21_PULLEN),
  .pullsel(`DP0_21_PULLSEL),
  .pad_pd(`DP0_21)
));
ap_DP0_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_21),
  .pullen(`DP0_21_PULLEN),
  .pullsel(`DP0_21_PULLSEL)
));
ap_DP0_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE)
));
ap_DP0_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_22_PINCTRL_0_IE),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_22),
  .pad(`DP0_22),
  .default_value(`default_value)));
ap_DP0_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE)
));
ap_DP0_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_22_PINCTRL_0_IE),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_22),
  .pad(`DP0_22),
  .default_value(`default_value)));
ap_DP0_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE)
));
ap_DP0_22_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_22_PINCTRL_0_IE),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_22),
  .pad(`DP0_22),
  .default_value(`default_value)));
ap_DP0_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_22_OUTFUNC_SEL),
  .gpioouten(`DP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`DP0_22_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`DP0_22),
  .pad_gz(`DP0_22_pad_y)
));
ap_DP0_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_22)
));
ap_DP0_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE)
));
ap_DP0_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_22_PINCTRL_0_IE),
  .outen(`DP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_22),
  .pad(`DP0_22),
  .default_value(`default_value)));
ap_DP0_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_22_PULLEN),
  .pullsel(`DP0_22_PULLSEL),
  .pad_pullup(`DP0_22)
));
ap_DP0_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .pullsel(`DP0_22_PULLSEL)
));
ap_DP0_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_22_PULLEN),
  .pullsel(`DP0_22_PULLSEL),
  .pad_pd(`DP0_22)
));
ap_DP0_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_22),
  .pullen(`DP0_22_PULLEN),
  .pullsel(`DP0_22_PULLSEL)
));
ap_DP0_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE)
));
ap_DP0_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_23_PINCTRL_0_IE),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_23),
  .pad(`DP0_23),
  .default_value(`default_value)));
ap_DP0_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE)
));
ap_DP0_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_23_PINCTRL_0_IE),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_23),
  .pad(`DP0_23),
  .default_value(`default_value)));
ap_DP0_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE)
));
ap_DP0_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_23_PINCTRL_0_IE),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_23),
  .pad(`DP0_23),
  .default_value(`default_value)));
ap_DP0_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE)
));
ap_DP0_23_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_23_PINCTRL_0_IE),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_23),
  .pad(`DP0_23),
  .default_value(`default_value)));
ap_DP0_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_23_OUTFUNC_SEL),
  .gpioouten(`DP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`DP0_23_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`DP0_23),
  .pad_gz(`DP0_23_pad_y)
));
ap_DP0_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_23)
));
ap_DP0_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE)
));
ap_DP0_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_23_PINCTRL_0_IE),
  .outen(`DP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_23),
  .pad(`DP0_23),
  .default_value(`default_value)));
ap_DP0_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_23_PULLEN),
  .pullsel(`DP0_23_PULLSEL),
  .pad_pullup(`DP0_23)
));
ap_DP0_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .pullsel(`DP0_23_PULLSEL)
));
ap_DP0_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_23_PULLEN),
  .pullsel(`DP0_23_PULLSEL),
  .pad_pd(`DP0_23)
));
ap_DP0_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_23),
  .pullen(`DP0_23_PULLEN),
  .pullsel(`DP0_23_PULLSEL)
));
ap_DP0_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE)
));
ap_DP0_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_24_PINCTRL_0_IE),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_24),
  .pad(`DP0_24),
  .default_value(`default_value)));
ap_DP0_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE)
));
ap_DP0_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_24_PINCTRL_0_IE),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_24),
  .pad(`DP0_24),
  .default_value(`default_value)));
ap_DP0_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE)
));
ap_DP0_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_24_PINCTRL_0_IE),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_24),
  .pad(`DP0_24),
  .default_value(`default_value)));
ap_DP0_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE)
));
ap_DP0_24_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_24_PINCTRL_0_IE),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_24),
  .pad(`DP0_24),
  .default_value(`default_value)));
ap_DP0_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_24_OUTFUNC_SEL),
  .gpioouten(`DP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`DP0_24_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`DP0_24),
  .pad_gz(`DP0_24_pad_y)
));
ap_DP0_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_24)
));
ap_DP0_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE)
));
ap_DP0_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_24_PINCTRL_0_IE),
  .outen(`DP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_24),
  .pad(`DP0_24),
  .default_value(`default_value)));
ap_DP0_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_24_PULLEN),
  .pullsel(`DP0_24_PULLSEL),
  .pad_pullup(`DP0_24)
));
ap_DP0_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .pullsel(`DP0_24_PULLSEL)
));
ap_DP0_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_24_PULLEN),
  .pullsel(`DP0_24_PULLSEL),
  .pad_pd(`DP0_24)
));
ap_DP0_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_24),
  .pullen(`DP0_24_PULLEN),
  .pullsel(`DP0_24_PULLSEL)
));
ap_DP0_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE)
));
ap_DP0_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_25_PINCTRL_0_IE),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_25),
  .pad(`DP0_25),
  .default_value(`default_value)));
ap_DP0_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE)
));
ap_DP0_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_25_PINCTRL_0_IE),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_25),
  .pad(`DP0_25),
  .default_value(`default_value)));
ap_DP0_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE)
));
ap_DP0_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_25_PINCTRL_0_IE),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_25),
  .pad(`DP0_25),
  .default_value(`default_value)));
ap_DP0_25_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE)
));
ap_DP0_25_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP0_25_PINCTRL_0_IE),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_25),
  .pad(`DP0_25),
  .default_value(`default_value)));
ap_DP0_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_25_OUTFUNC_SEL),
  .gpioouten(`DP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP0_25_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP0_25),
  .pad_gz(`DP0_25_pad_y)
));
ap_DP0_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_25)
));
ap_DP0_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE)
));
ap_DP0_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_25_PINCTRL_0_IE),
  .outen(`DP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_25),
  .pad(`DP0_25),
  .default_value(`default_value)));
ap_DP0_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_25_PULLEN),
  .pullsel(`DP0_25_PULLSEL),
  .pad_pullup(`DP0_25)
));
ap_DP0_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .pullsel(`DP0_25_PULLSEL)
));
ap_DP0_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_25_PULLEN),
  .pullsel(`DP0_25_PULLSEL),
  .pad_pd(`DP0_25)
));
ap_DP0_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_25),
  .pullen(`DP0_25_PULLEN),
  .pullsel(`DP0_25_PULLSEL)
));
ap_DP0_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE)
));
ap_DP0_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_26_PINCTRL_0_IE),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_26),
  .pad(`DP0_26),
  .default_value(`default_value)));
ap_DP0_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE)
));
ap_DP0_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_26_PINCTRL_0_IE),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_26),
  .pad(`DP0_26),
  .default_value(`default_value)));
ap_DP0_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE)
));
ap_DP0_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_26_PINCTRL_0_IE),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_26),
  .pad(`DP0_26),
  .default_value(`default_value)));
ap_DP0_26_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_26_OUTFUNC_SEL),
  .gpioouten(`DP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP0_26_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP0_26),
  .pad_gz(`DP0_26_pad_y)
));
ap_DP0_26_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_26)
));
ap_DP0_26_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE)
));
ap_DP0_26_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_26_PINCTRL_0_IE),
  .outen(`DP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_26),
  .pad(`DP0_26),
  .default_value(`default_value)));
ap_DP0_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_26_PULLEN),
  .pullsel(`DP0_26_PULLSEL),
  .pad_pullup(`DP0_26)
));
ap_DP0_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .pullsel(`DP0_26_PULLSEL)
));
ap_DP0_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_26_PULLEN),
  .pullsel(`DP0_26_PULLSEL),
  .pad_pd(`DP0_26)
));
ap_DP0_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_26),
  .pullen(`DP0_26_PULLEN),
  .pullsel(`DP0_26_PULLSEL)
));
ap_DP0_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE)
));
ap_DP0_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_27_PINCTRL_0_IE),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_27),
  .pad(`DP0_27),
  .default_value(`default_value)));
ap_DP0_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE)
));
ap_DP0_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_27_PINCTRL_0_IE),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_27),
  .pad(`DP0_27),
  .default_value(`default_value)));
ap_DP0_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE)
));
ap_DP0_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_27_PINCTRL_0_IE),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_27),
  .pad(`DP0_27),
  .default_value(`default_value)));
ap_DP0_27_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_27_OUTFUNC_SEL),
  .gpioouten(`DP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`DP0_27_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`DP0_27),
  .pad_gz(`DP0_27_pad_y)
));
ap_DP0_27_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_27)
));
ap_DP0_27_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE)
));
ap_DP0_27_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP0_27_PINCTRL_0_IE),
  .outen(`DP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_27),
  .pad(`DP0_27),
  .default_value(`default_value)));
ap_DP0_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_27_PULLEN),
  .pullsel(`DP0_27_PULLSEL),
  .pad_pullup(`DP0_27)
));
ap_DP0_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .pullsel(`DP0_27_PULLSEL)
));
ap_DP0_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_27_PULLEN),
  .pullsel(`DP0_27_PULLSEL),
  .pad_pd(`DP0_27)
));
ap_DP0_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_27),
  .pullen(`DP0_27_PULLEN),
  .pullsel(`DP0_27_PULLSEL)
));
ap_DP0_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`DP0_28),
  .pad_gz(`DP0_28_pad_y)
));
ap_DP0_28_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_28),
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE)
));
ap_DP0_28_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_28_PINCTRL_0_IE),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_28),
  .pad(`DP0_28),
  .default_value(`default_value)));
ap_DP0_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP0_28),
  .pad_gz(`DP0_28_pad_y)
));
ap_DP0_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_28),
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE)
));
ap_DP0_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_28_PINCTRL_0_IE),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_28),
  .pad(`DP0_28),
  .default_value(`default_value)));
ap_DP0_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP0_28),
  .pad_gz(`DP0_28_pad_y)
));
ap_DP0_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXCLK_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`FSI2RXCLK_OUT),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXCLK_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`FSI2RXCLK_OUT),
  .pad(`DP0_28),
  .pad_gz(`DP0_28_pad_y)
));
ap_DP0_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_28),
  .pullen(`DP0_28_PULLEN),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE)
));
ap_DP0_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_28_PINCTRL_0_IE),
  .outen(`DP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_28),
  .pad(`DP0_28),
  .default_value(`default_value)));
ap_DP0_28_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP0_28)
));
ap_DP0_28_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_28_OUTFUNC_SEL),
  .gpioouten(`DP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP0_28_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP0_28),
  .pad_gz(`DP0_28_pad_y)
));
ap_DP0_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_28_PULLEN),
  .pullsel(`DP0_28_PULLSEL),
  .pad_pullup(`DP0_28)
));
ap_DP0_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_28),
  .pullen(`DP0_28_PULLEN),
  .pullsel(`DP0_28_PULLSEL)
));
ap_DP0_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_28_PULLEN),
  .pullsel(`DP0_28_PULLSEL),
  .pad_pd(`DP0_28)
));
ap_DP0_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_28),
  .pullen(`DP0_28_PULLEN),
  .pullsel(`DP0_28_PULLSEL)
));
ap_DP0_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`DP0_29),
  .pad_gz(`DP0_29_pad_y)
));
ap_DP0_29_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_29),
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE)
));
ap_DP0_29_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_29_PINCTRL_0_IE),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_29),
  .pad(`DP0_29),
  .default_value(`default_value)));
ap_DP0_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP0_29),
  .pad_gz(`DP0_29_pad_y)
));
ap_DP0_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_29),
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE)
));
ap_DP0_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_29_PINCTRL_0_IE),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_29),
  .pad(`DP0_29),
  .default_value(`default_value)));
ap_DP0_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP0_29),
  .pad_gz(`DP0_29_pad_y)
));
ap_DP0_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD0_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`FSI2RXD0_OUT),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD0_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`FSI2RXD0_OUT),
  .pad(`DP0_29),
  .pad_gz(`DP0_29_pad_y)
));
ap_DP0_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_29),
  .pullen(`DP0_29_PULLEN),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE)
));
ap_DP0_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_29_PINCTRL_0_IE),
  .outen(`DP0_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_29),
  .pad(`DP0_29),
  .default_value(`default_value)));
ap_DP0_29_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP0_29)
));
ap_DP0_29_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_29_OUTFUNC_SEL),
  .gpioouten(`DP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP0_29_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP0_29),
  .pad_gz(`DP0_29_pad_y)
));
ap_DP0_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_29_PULLEN),
  .pullsel(`DP0_29_PULLSEL),
  .pad_pullup(`DP0_29)
));
ap_DP0_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_29),
  .pullen(`DP0_29_PULLEN),
  .pullsel(`DP0_29_PULLSEL)
));
ap_DP0_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_29_PULLEN),
  .pullsel(`DP0_29_PULLSEL),
  .pad_pd(`DP0_29)
));
ap_DP0_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_29),
  .pullen(`DP0_29_PULLEN),
  .pullsel(`DP0_29_PULLSEL)
));
ap_DP0_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`DP0_30),
  .pad_gz(`DP0_30_pad_y)
));
ap_DP0_30_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_30),
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE)
));
ap_DP0_30_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_30_PINCTRL_0_IE),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_30),
  .pad(`DP0_30),
  .default_value(`default_value)));
ap_DP0_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP0_30),
  .pad_gz(`DP0_30_pad_y)
));
ap_DP0_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_30),
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE)
));
ap_DP0_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_30_PINCTRL_0_IE),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_30),
  .pad(`DP0_30),
  .default_value(`default_value)));
ap_DP0_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP0_30),
  .pad_gz(`DP0_30_pad_y)
));
ap_DP0_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD1_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`FSI2RXD1_OUT),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD1_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`FSI2RXD1_OUT),
  .pad(`DP0_30),
  .pad_gz(`DP0_30_pad_y)
));
ap_DP0_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_30),
  .pullen(`DP0_30_PULLEN),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE)
));
ap_DP0_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_30_PINCTRL_0_IE),
  .outen(`DP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_30),
  .pad(`DP0_30),
  .default_value(`default_value)));
ap_DP0_30_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP0_30)
));
ap_DP0_30_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_30_OUTFUNC_SEL),
  .gpioouten(`DP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP0_30_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP0_30),
  .pad_gz(`DP0_30_pad_y)
));
ap_DP0_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_30_PULLEN),
  .pullsel(`DP0_30_PULLSEL),
  .pad_pullup(`DP0_30)
));
ap_DP0_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_30),
  .pullen(`DP0_30_PULLEN),
  .pullsel(`DP0_30_PULLSEL)
));
ap_DP0_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_30_PULLEN),
  .pullsel(`DP0_30_PULLSEL),
  .pad_pd(`DP0_30)
));
ap_DP0_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_30),
  .pullen(`DP0_30_PULLEN),
  .pullsel(`DP0_30_PULLSEL)
));
ap_DP0_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`DP0_31),
  .pad_gz(`DP0_31_pad_y)
));
ap_DP0_31_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_31),
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE)
));
ap_DP0_31_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP0_31_PINCTRL_0_IE),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_31),
  .pad(`DP0_31),
  .default_value(`default_value)));
ap_DP0_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP0_31),
  .pad_gz(`DP0_31_pad_y)
));
ap_DP0_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_31),
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE)
));
ap_DP0_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP0_31_PINCTRL_0_IE),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_31),
  .pad(`DP0_31),
  .default_value(`default_value)));
ap_DP0_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP0_31),
  .pad_gz(`DP0_31_pad_y)
));
ap_DP0_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXCLK_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`FSI3TXCLK_OUT),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXCLK_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`FSI3TXCLK_OUT),
  .pad(`DP0_31),
  .pad_gz(`DP0_31_pad_y)
));
ap_DP0_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP0_31),
  .pullen(`DP0_31_PULLEN),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE)
));
ap_DP0_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP0_31_PINCTRL_0_IE),
  .outen(`DP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP0_31),
  .pad(`DP0_31),
  .default_value(`default_value)));
ap_DP0_31_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP0_31)
));
ap_DP0_31_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP0_31_OUTFUNC_SEL),
  .gpioouten(`DP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP0_31_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP0_31),
  .pad_gz(`DP0_31_pad_y)
));
ap_DP0_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP0_31_PULLEN),
  .pullsel(`DP0_31_PULLSEL),
  .pad_pullup(`DP0_31)
));
ap_DP0_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP0_31),
  .pullen(`DP0_31_PULLEN),
  .pullsel(`DP0_31_PULLSEL)
));
ap_DP0_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP0_31_PULLEN),
  .pullsel(`DP0_31_PULLSEL),
  .pad_pd(`DP0_31)
));
ap_DP0_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP0_31),
  .pullen(`DP0_31_PULLEN),
  .pullsel(`DP0_31_PULLSEL)
));
ap_DP1_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP1_0),
  .pad_gz(`DP1_0_pad_y)
));
ap_DP1_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP1_0),
  .pad_gz(`DP1_0_pad_y)
));
ap_DP1_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_0_PULLEN),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_0),
  .pullen(`DP1_0_PULLEN),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE)
));
ap_DP1_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_0_PINCTRL_0_IE),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_0),
  .pad(`DP1_0),
  .default_value(`default_value)));
ap_DP1_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP1_0),
  .pad_gz(`DP1_0_pad_y)
));
ap_DP1_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_0_PULLEN),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_0),
  .pullen(`DP1_0_PULLEN),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE)
));
ap_DP1_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_0_PINCTRL_0_IE),
  .outen(`DP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_0),
  .pad(`DP1_0),
  .default_value(`default_value)));
ap_DP1_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP1_0)
));
ap_DP1_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_0_OUTFUNC_SEL),
  .gpioouten(`DP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP1_0_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP1_0),
  .pad_gz(`DP1_0_pad_y)
));
ap_DP1_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_0_PULLEN),
  .pullsel(`DP1_0_PULLSEL),
  .pad_pullup(`DP1_0)
));
ap_DP1_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_0),
  .pullen(`DP1_0_PULLEN),
  .pullsel(`DP1_0_PULLSEL)
));
ap_DP1_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_0_PULLEN),
  .pullsel(`DP1_0_PULLSEL),
  .pad_pd(`DP1_0)
));
ap_DP1_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_0),
  .pullen(`DP1_0_PULLEN),
  .pullsel(`DP1_0_PULLSEL)
));
ap_DP1_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP1_1),
  .pad_gz(`DP1_1_pad_y)
));
ap_DP1_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP1_1),
  .pad_gz(`DP1_1_pad_y)
));
ap_DP1_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_1_PULLEN),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_1),
  .pullen(`DP1_1_PULLEN),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE)
));
ap_DP1_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_1_PINCTRL_0_IE),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_1),
  .pad(`DP1_1),
  .default_value(`default_value)));
ap_DP1_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP1_1),
  .pad_gz(`DP1_1_pad_y)
));
ap_DP1_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_1_PULLEN),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_1),
  .pullen(`DP1_1_PULLEN),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE)
));
ap_DP1_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_1_PINCTRL_0_IE),
  .outen(`DP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_1),
  .pad(`DP1_1),
  .default_value(`default_value)));
ap_DP1_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP1_1)
));
ap_DP1_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_1_OUTFUNC_SEL),
  .gpioouten(`DP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP1_1_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP1_1),
  .pad_gz(`DP1_1_pad_y)
));
ap_DP1_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_1_PULLEN),
  .pullsel(`DP1_1_PULLSEL),
  .pad_pullup(`DP1_1)
));
ap_DP1_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_1),
  .pullen(`DP1_1_PULLEN),
  .pullsel(`DP1_1_PULLSEL)
));
ap_DP1_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_1_PULLEN),
  .pullsel(`DP1_1_PULLSEL),
  .pad_pd(`DP1_1)
));
ap_DP1_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_1),
  .pullen(`DP1_1_PULLEN),
  .pullsel(`DP1_1_PULLSEL)
));
ap_DP1_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP1_2),
  .pad_gz(`DP1_2_pad_y)
));
ap_DP1_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP1_2),
  .pad_gz(`DP1_2_pad_y)
));
ap_DP1_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_2_PULLEN),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_2),
  .pullen(`DP1_2_PULLEN),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE)
));
ap_DP1_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_2_PINCTRL_0_IE),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_2),
  .pad(`DP1_2),
  .default_value(`default_value)));
ap_DP1_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP1_2),
  .pad_gz(`DP1_2_pad_y)
));
ap_DP1_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_2_PULLEN),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_2),
  .pullen(`DP1_2_PULLEN),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE)
));
ap_DP1_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_2_PINCTRL_0_IE),
  .outen(`DP1_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_2),
  .pad(`DP1_2),
  .default_value(`default_value)));
ap_DP1_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP1_2)
));
ap_DP1_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_2_OUTFUNC_SEL),
  .gpioouten(`DP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP1_2_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP1_2),
  .pad_gz(`DP1_2_pad_y)
));
ap_DP1_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_2_PULLEN),
  .pullsel(`DP1_2_PULLSEL),
  .pad_pullup(`DP1_2)
));
ap_DP1_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_2),
  .pullen(`DP1_2_PULLEN),
  .pullsel(`DP1_2_PULLSEL)
));
ap_DP1_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_2_PULLEN),
  .pullsel(`DP1_2_PULLSEL),
  .pad_pd(`DP1_2)
));
ap_DP1_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_2),
  .pullen(`DP1_2_PULLEN),
  .pullsel(`DP1_2_PULLSEL)
));
ap_DP1_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP1_3),
  .pad_gz(`DP1_3_pad_y)
));
ap_DP1_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP1_3),
  .pad_gz(`DP1_3_pad_y)
));
ap_DP1_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_3_PULLEN),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_3),
  .pullen(`DP1_3_PULLEN),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE)
));
ap_DP1_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_3_PINCTRL_0_IE),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_3),
  .pad(`DP1_3),
  .default_value(`default_value)));
ap_DP1_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP1_3),
  .pad_gz(`DP1_3_pad_y)
));
ap_DP1_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_3_PULLEN),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_3),
  .pullen(`DP1_3_PULLEN),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE)
));
ap_DP1_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_3_PINCTRL_0_IE),
  .outen(`DP1_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_3),
  .pad(`DP1_3),
  .default_value(`default_value)));
ap_DP1_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP1_3)
));
ap_DP1_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_3_OUTFUNC_SEL),
  .gpioouten(`DP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP1_3_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP1_3),
  .pad_gz(`DP1_3_pad_y)
));
ap_DP1_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_3_PULLEN),
  .pullsel(`DP1_3_PULLSEL),
  .pad_pullup(`DP1_3)
));
ap_DP1_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_3),
  .pullen(`DP1_3_PULLEN),
  .pullsel(`DP1_3_PULLSEL)
));
ap_DP1_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_3_PULLEN),
  .pullsel(`DP1_3_PULLSEL),
  .pad_pd(`DP1_3)
));
ap_DP1_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_3),
  .pullen(`DP1_3_PULLEN),
  .pullsel(`DP1_3_PULLSEL)
));
ap_DP1_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP1_4),
  .pad_gz(`DP1_4_pad_y)
));
ap_DP1_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP1_4),
  .pad_gz(`DP1_4_pad_y)
));
ap_DP1_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_4_PULLEN),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_4),
  .pullen(`DP1_4_PULLEN),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE)
));
ap_DP1_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_4_PINCTRL_0_IE),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_4),
  .pad(`DP1_4),
  .default_value(`default_value)));
ap_DP1_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP1_4),
  .pad_gz(`DP1_4_pad_y)
));
ap_DP1_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_4_PULLEN),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_4),
  .pullen(`DP1_4_PULLEN),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE)
));
ap_DP1_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_4_PINCTRL_0_IE),
  .outen(`DP1_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_4),
  .pad(`DP1_4),
  .default_value(`default_value)));
ap_DP1_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP1_4)
));
ap_DP1_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_4_OUTFUNC_SEL),
  .gpioouten(`DP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP1_4_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP1_4),
  .pad_gz(`DP1_4_pad_y)
));
ap_DP1_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_4_PULLEN),
  .pullsel(`DP1_4_PULLSEL),
  .pad_pullup(`DP1_4)
));
ap_DP1_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_4),
  .pullen(`DP1_4_PULLEN),
  .pullsel(`DP1_4_PULLSEL)
));
ap_DP1_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_4_PULLEN),
  .pullsel(`DP1_4_PULLSEL),
  .pad_pd(`DP1_4)
));
ap_DP1_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_4),
  .pullen(`DP1_4_PULLEN),
  .pullsel(`DP1_4_PULLSEL)
));
ap_DP1_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP1_5),
  .pad_gz(`DP1_5_pad_y)
));
ap_DP1_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP1_5),
  .pad_gz(`DP1_5_pad_y)
));
ap_DP1_5_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_5_PULLEN),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_5),
  .pullen(`DP1_5_PULLEN),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE)
));
ap_DP1_5_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_5_PINCTRL_0_IE),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_5),
  .pad(`DP1_5),
  .default_value(`default_value)));
ap_DP1_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP1_5),
  .pad_gz(`DP1_5_pad_y)
));
ap_DP1_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_5_PULLEN),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_5),
  .pullen(`DP1_5_PULLEN),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE)
));
ap_DP1_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_5_PINCTRL_0_IE),
  .outen(`DP1_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_5),
  .pad(`DP1_5),
  .default_value(`default_value)));
ap_DP1_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP1_5)
));
ap_DP1_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_5_OUTFUNC_SEL),
  .gpioouten(`DP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP1_5_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP1_5),
  .pad_gz(`DP1_5_pad_y)
));
ap_DP1_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_5_PULLEN),
  .pullsel(`DP1_5_PULLSEL),
  .pad_pullup(`DP1_5)
));
ap_DP1_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_5),
  .pullen(`DP1_5_PULLEN),
  .pullsel(`DP1_5_PULLSEL)
));
ap_DP1_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_5_PULLEN),
  .pullsel(`DP1_5_PULLSEL),
  .pad_pd(`DP1_5)
));
ap_DP1_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_5),
  .pullen(`DP1_5_PULLEN),
  .pullsel(`DP1_5_PULLSEL)
));
ap_DP1_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP1_6),
  .pad_gz(`DP1_6_pad_y)
));
ap_DP1_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP1_6),
  .pad_gz(`DP1_6_pad_y)
));
ap_DP1_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_6_PULLEN),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_6),
  .pullen(`DP1_6_PULLEN),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE)
));
ap_DP1_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_6_PINCTRL_0_IE),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_6),
  .pad(`DP1_6),
  .default_value(`default_value)));
ap_DP1_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP1_6),
  .pad_gz(`DP1_6_pad_y)
));
ap_DP1_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_6_PULLEN),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_6),
  .pullen(`DP1_6_PULLEN),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE)
));
ap_DP1_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_6_PINCTRL_0_IE),
  .outen(`DP1_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_6),
  .pad(`DP1_6),
  .default_value(`default_value)));
ap_DP1_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP1_6)
));
ap_DP1_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_6_OUTFUNC_SEL),
  .gpioouten(`DP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP1_6_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP1_6),
  .pad_gz(`DP1_6_pad_y)
));
ap_DP1_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_6_PULLEN),
  .pullsel(`DP1_6_PULLSEL),
  .pad_pullup(`DP1_6)
));
ap_DP1_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_6),
  .pullen(`DP1_6_PULLEN),
  .pullsel(`DP1_6_PULLSEL)
));
ap_DP1_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_6_PULLEN),
  .pullsel(`DP1_6_PULLSEL),
  .pad_pd(`DP1_6)
));
ap_DP1_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_6),
  .pullen(`DP1_6_PULLEN),
  .pullsel(`DP1_6_PULLSEL)
));
ap_DP1_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP1_7),
  .pad_gz(`DP1_7_pad_y)
));
ap_DP1_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP1_7),
  .pad_gz(`DP1_7_pad_y)
));
ap_DP1_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_7_PULLEN),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_7),
  .pullen(`DP1_7_PULLEN),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE)
));
ap_DP1_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_7_PINCTRL_0_IE),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_7),
  .pad(`DP1_7),
  .default_value(`default_value)));
ap_DP1_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP1_7),
  .pad_gz(`DP1_7_pad_y)
));
ap_DP1_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_7_PULLEN),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_7),
  .pullen(`DP1_7_PULLEN),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE)
));
ap_DP1_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_7_PINCTRL_0_IE),
  .outen(`DP1_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_7),
  .pad(`DP1_7),
  .default_value(`default_value)));
ap_DP1_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP1_7)
));
ap_DP1_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_7_OUTFUNC_SEL),
  .gpioouten(`DP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP1_7_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP1_7),
  .pad_gz(`DP1_7_pad_y)
));
ap_DP1_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_7_PULLEN),
  .pullsel(`DP1_7_PULLSEL),
  .pad_pullup(`DP1_7)
));
ap_DP1_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_7),
  .pullen(`DP1_7_PULLEN),
  .pullsel(`DP1_7_PULLSEL)
));
ap_DP1_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_7_PULLEN),
  .pullsel(`DP1_7_PULLSEL),
  .pad_pd(`DP1_7)
));
ap_DP1_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_7),
  .pullen(`DP1_7_PULLEN),
  .pullsel(`DP1_7_PULLSEL)
));
ap_DP1_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP1_8)
));
ap_DP1_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP1_8),
  .pad_gz(`DP1_8_pad_y)
));
ap_DP1_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP1_8)
));
ap_DP1_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP1_8),
  .pad_gz(`DP1_8_pad_y)
));
ap_DP1_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_8_PULLEN),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_8)
));
ap_DP1_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_8),
  .pullen(`DP1_8_PULLEN),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE)
));
ap_DP1_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_8_PINCTRL_0_IE),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_8),
  .pad(`DP1_8),
  .default_value(`default_value)));
ap_DP1_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP1_8)
));
ap_DP1_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_8_OUTFUNC_SEL),
  .gpioouten(`DP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP1_8_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP1_8),
  .pad_gz(`DP1_8_pad_y)
));
ap_DP1_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_8_PULLEN),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_8)
));
ap_DP1_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_8),
  .pullen(`DP1_8_PULLEN),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE)
));
ap_DP1_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_8_PINCTRL_0_IE),
  .outen(`DP1_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_8),
  .pad(`DP1_8),
  .default_value(`default_value)));
ap_DP1_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_8_PULLEN),
  .pullsel(`DP1_8_PULLSEL),
  .pad_pullup(`DP1_8)
));
ap_DP1_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_8),
  .pullen(`DP1_8_PULLEN),
  .pullsel(`DP1_8_PULLSEL)
));
ap_DP1_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_8_PULLEN),
  .pullsel(`DP1_8_PULLSEL),
  .pad_pd(`DP1_8)
));
ap_DP1_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_8),
  .pullen(`DP1_8_PULLEN),
  .pullsel(`DP1_8_PULLSEL)
));
ap_DP1_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP1_9)
));
ap_DP1_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP1_9),
  .pad_gz(`DP1_9_pad_y)
));
ap_DP1_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP1_9)
));
ap_DP1_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP1_9),
  .pad_gz(`DP1_9_pad_y)
));
ap_DP1_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_9_PULLEN),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_9)
));
ap_DP1_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_9),
  .pullen(`DP1_9_PULLEN),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE)
));
ap_DP1_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_9_PINCTRL_0_IE),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_9),
  .pad(`DP1_9),
  .default_value(`default_value)));
ap_DP1_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP1_9)
));
ap_DP1_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_9_OUTFUNC_SEL),
  .gpioouten(`DP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP1_9_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP1_9),
  .pad_gz(`DP1_9_pad_y)
));
ap_DP1_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_9_PULLEN),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_9)
));
ap_DP1_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_9),
  .pullen(`DP1_9_PULLEN),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE)
));
ap_DP1_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_9_PINCTRL_0_IE),
  .outen(`DP1_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_9),
  .pad(`DP1_9),
  .default_value(`default_value)));
ap_DP1_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_9_PULLEN),
  .pullsel(`DP1_9_PULLSEL),
  .pad_pullup(`DP1_9)
));
ap_DP1_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_9),
  .pullen(`DP1_9_PULLEN),
  .pullsel(`DP1_9_PULLSEL)
));
ap_DP1_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_9_PULLEN),
  .pullsel(`DP1_9_PULLSEL),
  .pad_pd(`DP1_9)
));
ap_DP1_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_9),
  .pullen(`DP1_9_PULLEN),
  .pullsel(`DP1_9_PULLSEL)
));
ap_DP1_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_10_OUTFUNC_SEL),
  .gpioouten(`DP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP1_10_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP1_10)
));
ap_DP1_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_10_OUTFUNC_SEL),
  .gpioouten(`DP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP1_10_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP1_10),
  .pad_gz(`DP1_10_pad_y)
));
ap_DP1_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_10_OUTFUNC_SEL),
  .gpioouten(`DP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP1_10_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP1_10)
));
ap_DP1_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_10_OUTFUNC_SEL),
  .gpioouten(`DP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP1_10_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP1_10),
  .pad_gz(`DP1_10_pad_y)
));
ap_DP1_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_10_PULLEN),
  .outen(`DP1_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_10)
));
ap_DP1_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_10),
  .pullen(`DP1_10_PULLEN),
  .outen(`DP1_10_GPIO_OUTPUT_ENABLE)
));
ap_DP1_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_10_PINCTRL_0_IE),
  .outen(`DP1_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_10),
  .pad(`DP1_10),
  .default_value(`default_value)));
ap_DP1_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_10_PULLEN),
  .pullsel(`DP1_10_PULLSEL),
  .pad_pullup(`DP1_10)
));
ap_DP1_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_10),
  .pullen(`DP1_10_PULLEN),
  .pullsel(`DP1_10_PULLSEL)
));
ap_DP1_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_10_PULLEN),
  .pullsel(`DP1_10_PULLSEL),
  .pad_pd(`DP1_10)
));
ap_DP1_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_10),
  .pullen(`DP1_10_PULLEN),
  .pullsel(`DP1_10_PULLSEL)
));
ap_DP1_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_11_OUTFUNC_SEL),
  .gpioouten(`DP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP1_11_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP1_11)
));
ap_DP1_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_11_OUTFUNC_SEL),
  .gpioouten(`DP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP1_11_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP1_11),
  .pad_gz(`DP1_11_pad_y)
));
ap_DP1_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_11_OUTFUNC_SEL),
  .gpioouten(`DP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP1_11_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP1_11)
));
ap_DP1_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_11_OUTFUNC_SEL),
  .gpioouten(`DP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP1_11_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP1_11),
  .pad_gz(`DP1_11_pad_y)
));
ap_DP1_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_11_PULLEN),
  .outen(`DP1_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_11)
));
ap_DP1_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_11),
  .pullen(`DP1_11_PULLEN),
  .outen(`DP1_11_GPIO_OUTPUT_ENABLE)
));
ap_DP1_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_11_PINCTRL_0_IE),
  .outen(`DP1_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_11),
  .pad(`DP1_11),
  .default_value(`default_value)));
ap_DP1_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_11_PULLEN),
  .pullsel(`DP1_11_PULLSEL),
  .pad_pullup(`DP1_11)
));
ap_DP1_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_11),
  .pullen(`DP1_11_PULLEN),
  .pullsel(`DP1_11_PULLSEL)
));
ap_DP1_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_11_PULLEN),
  .pullsel(`DP1_11_PULLSEL),
  .pad_pd(`DP1_11)
));
ap_DP1_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_11),
  .pullen(`DP1_11_PULLEN),
  .pullsel(`DP1_11_PULLSEL)
));
ap_DP1_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_12_OUTFUNC_SEL),
  .gpioouten(`DP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP1_12_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP1_12)
));
ap_DP1_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_12_OUTFUNC_SEL),
  .gpioouten(`DP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP1_12_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP1_12),
  .pad_gz(`DP1_12_pad_y)
));
ap_DP1_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_12_OUTFUNC_SEL),
  .gpioouten(`DP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP1_12_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP1_12)
));
ap_DP1_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_12_OUTFUNC_SEL),
  .gpioouten(`DP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP1_12_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP1_12),
  .pad_gz(`DP1_12_pad_y)
));
ap_DP1_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_12_PULLEN),
  .outen(`DP1_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_12)
));
ap_DP1_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_12),
  .pullen(`DP1_12_PULLEN),
  .outen(`DP1_12_GPIO_OUTPUT_ENABLE)
));
ap_DP1_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_12_PINCTRL_0_IE),
  .outen(`DP1_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_12),
  .pad(`DP1_12),
  .default_value(`default_value)));
ap_DP1_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_12_PULLEN),
  .pullsel(`DP1_12_PULLSEL),
  .pad_pullup(`DP1_12)
));
ap_DP1_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_12),
  .pullen(`DP1_12_PULLEN),
  .pullsel(`DP1_12_PULLSEL)
));
ap_DP1_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_12_PULLEN),
  .pullsel(`DP1_12_PULLSEL),
  .pad_pd(`DP1_12)
));
ap_DP1_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_12),
  .pullen(`DP1_12_PULLEN),
  .pullsel(`DP1_12_PULLSEL)
));
ap_DP1_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP1_13),
  .pad_gz(`DP1_13_pad_y)
));
ap_DP1_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP1_13),
  .pad_gz(`DP1_13_pad_y)
));
ap_DP1_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_13),
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE)
));
ap_DP1_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_13_PINCTRL_0_IE),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_13),
  .pad(`DP1_13),
  .default_value(`default_value)));
ap_DP1_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`DP1_13),
  .pad_gz(`DP1_13_pad_y)
));
ap_DP1_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_13),
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE)
));
ap_DP1_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_13_PINCTRL_0_IE),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_13),
  .pad(`DP1_13),
  .default_value(`default_value)));
ap_DP1_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_13_OUTFUNC_SEL),
  .gpioouten(`DP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`DP1_13_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`DP1_13),
  .pad_gz(`DP1_13_pad_y)
));
ap_DP1_13_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_13)
));
ap_DP1_13_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_13),
  .pullen(`DP1_13_PULLEN),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE)
));
ap_DP1_13_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_13_PINCTRL_0_IE),
  .outen(`DP1_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_13),
  .pad(`DP1_13),
  .default_value(`default_value)));
ap_DP1_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_13_PULLEN),
  .pullsel(`DP1_13_PULLSEL),
  .pad_pullup(`DP1_13)
));
ap_DP1_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_13),
  .pullen(`DP1_13_PULLEN),
  .pullsel(`DP1_13_PULLSEL)
));
ap_DP1_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_13_PULLEN),
  .pullsel(`DP1_13_PULLSEL),
  .pad_pd(`DP1_13)
));
ap_DP1_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_13),
  .pullen(`DP1_13_PULLEN),
  .pullsel(`DP1_13_PULLSEL)
));
ap_DP1_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP1_14),
  .pad_gz(`DP1_14_pad_y)
));
ap_DP1_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP1_14),
  .pad_gz(`DP1_14_pad_y)
));
ap_DP1_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_14),
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE)
));
ap_DP1_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_14_PINCTRL_0_IE),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_14),
  .pad(`DP1_14),
  .default_value(`default_value)));
ap_DP1_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`DP1_14),
  .pad_gz(`DP1_14_pad_y)
));
ap_DP1_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_14),
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE)
));
ap_DP1_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_14_PINCTRL_0_IE),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_14),
  .pad(`DP1_14),
  .default_value(`default_value)));
ap_DP1_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_14_OUTFUNC_SEL),
  .gpioouten(`DP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`DP1_14_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`DP1_14),
  .pad_gz(`DP1_14_pad_y)
));
ap_DP1_14_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_14)
));
ap_DP1_14_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_14),
  .pullen(`DP1_14_PULLEN),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE)
));
ap_DP1_14_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_14_PINCTRL_0_IE),
  .outen(`DP1_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_14),
  .pad(`DP1_14),
  .default_value(`default_value)));
ap_DP1_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_14_PULLEN),
  .pullsel(`DP1_14_PULLSEL),
  .pad_pullup(`DP1_14)
));
ap_DP1_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_14),
  .pullen(`DP1_14_PULLEN),
  .pullsel(`DP1_14_PULLSEL)
));
ap_DP1_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_14_PULLEN),
  .pullsel(`DP1_14_PULLSEL),
  .pad_pd(`DP1_14)
));
ap_DP1_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_14),
  .pullen(`DP1_14_PULLEN),
  .pullsel(`DP1_14_PULLSEL)
));
ap_DP1_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP1_15),
  .pad_gz(`DP1_15_pad_y)
));
ap_DP1_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP1_15),
  .pad_gz(`DP1_15_pad_y)
));
ap_DP1_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_15),
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE)
));
ap_DP1_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_15_PINCTRL_0_IE),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_15),
  .pad(`DP1_15),
  .default_value(`default_value)));
ap_DP1_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP1_15),
  .pad_gz(`DP1_15_pad_y)
));
ap_DP1_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_15),
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE)
));
ap_DP1_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_15_PINCTRL_0_IE),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_15),
  .pad(`DP1_15),
  .default_value(`default_value)));
ap_DP1_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_15_OUTFUNC_SEL),
  .gpioouten(`DP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`DP1_15_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`DP1_15),
  .pad_gz(`DP1_15_pad_y)
));
ap_DP1_15_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_15)
));
ap_DP1_15_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_15),
  .pullen(`DP1_15_PULLEN),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE)
));
ap_DP1_15_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_15_PINCTRL_0_IE),
  .outen(`DP1_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_15),
  .pad(`DP1_15),
  .default_value(`default_value)));
ap_DP1_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_15_PULLEN),
  .pullsel(`DP1_15_PULLSEL),
  .pad_pullup(`DP1_15)
));
ap_DP1_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_15),
  .pullen(`DP1_15_PULLEN),
  .pullsel(`DP1_15_PULLSEL)
));
ap_DP1_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_15_PULLEN),
  .pullsel(`DP1_15_PULLSEL),
  .pad_pd(`DP1_15)
));
ap_DP1_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_15),
  .pullen(`DP1_15_PULLEN),
  .pullsel(`DP1_15_PULLSEL)
));
ap_DP1_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP1_16),
  .pad_gz(`DP1_16_pad_y)
));
ap_DP1_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR0_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR0_OUT),
  .pad(`DP1_16),
  .pad_gz(`DP1_16_pad_y)
));
ap_DP1_16_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_16),
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE)
));
ap_DP1_16_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_16_PINCTRL_0_IE),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_16),
  .pad(`DP1_16),
  .default_value(`default_value)));
ap_DP1_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP1_16),
  .pad_gz(`DP1_16_pad_y)
));
ap_DP1_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_16),
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE)
));
ap_DP1_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_16_PINCTRL_0_IE),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_16),
  .pad(`DP1_16),
  .default_value(`default_value)));
ap_DP1_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_16_OUTFUNC_SEL),
  .gpioouten(`DP1_16_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`DP1_16_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`DP1_16),
  .pad_gz(`DP1_16_pad_y)
));
ap_DP1_16_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_16)
));
ap_DP1_16_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_16),
  .pullen(`DP1_16_PULLEN),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE)
));
ap_DP1_16_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_16_PINCTRL_0_IE),
  .outen(`DP1_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_16),
  .pad(`DP1_16),
  .default_value(`default_value)));
ap_DP1_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_16_PULLEN),
  .pullsel(`DP1_16_PULLSEL),
  .pad_pullup(`DP1_16)
));
ap_DP1_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_16),
  .pullen(`DP1_16_PULLEN),
  .pullsel(`DP1_16_PULLSEL)
));
ap_DP1_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_16_PULLEN),
  .pullsel(`DP1_16_PULLSEL),
  .pad_pd(`DP1_16)
));
ap_DP1_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_16),
  .pullen(`DP1_16_PULLEN),
  .pullsel(`DP1_16_PULLSEL)
));
ap_DP1_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP1_17),
  .pad_gz(`DP1_17_pad_y)
));
ap_DP1_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR1_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR1_OUT),
  .pad(`DP1_17),
  .pad_gz(`DP1_17_pad_y)
));
ap_DP1_17_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_17),
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE)
));
ap_DP1_17_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_17_PINCTRL_0_IE),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_17),
  .pad(`DP1_17),
  .default_value(`default_value)));
ap_DP1_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP1_17),
  .pad_gz(`DP1_17_pad_y)
));
ap_DP1_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_17),
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE)
));
ap_DP1_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_17_PINCTRL_0_IE),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_17),
  .pad(`DP1_17),
  .default_value(`default_value)));
ap_DP1_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_17_OUTFUNC_SEL),
  .gpioouten(`DP1_17_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`DP1_17_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`DP1_17),
  .pad_gz(`DP1_17_pad_y)
));
ap_DP1_17_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_17)
));
ap_DP1_17_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_17),
  .pullen(`DP1_17_PULLEN),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE)
));
ap_DP1_17_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_17_PINCTRL_0_IE),
  .outen(`DP1_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_17),
  .pad(`DP1_17),
  .default_value(`default_value)));
ap_DP1_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_17_PULLEN),
  .pullsel(`DP1_17_PULLSEL),
  .pad_pullup(`DP1_17)
));
ap_DP1_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_17),
  .pullen(`DP1_17_PULLEN),
  .pullsel(`DP1_17_PULLSEL)
));
ap_DP1_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_17_PULLEN),
  .pullsel(`DP1_17_PULLSEL),
  .pad_pd(`DP1_17)
));
ap_DP1_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_17),
  .pullen(`DP1_17_PULLEN),
  .pullsel(`DP1_17_PULLSEL)
));
ap_DP1_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP1_18),
  .pad_gz(`DP1_18_pad_y)
));
ap_DP1_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP1_18),
  .pad_gz(`DP1_18_pad_y)
));
ap_DP1_18_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_18),
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE)
));
ap_DP1_18_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_18_PINCTRL_0_IE),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_18),
  .pad(`DP1_18),
  .default_value(`default_value)));
ap_DP1_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP1_18),
  .pad_gz(`DP1_18_pad_y)
));
ap_DP1_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_18),
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE)
));
ap_DP1_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_18_PINCTRL_0_IE),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_18),
  .pad(`DP1_18),
  .default_value(`default_value)));
ap_DP1_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_18_OUTFUNC_SEL),
  .gpioouten(`DP1_18_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`DP1_18_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`DP1_18),
  .pad_gz(`DP1_18_pad_y)
));
ap_DP1_18_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_18)
));
ap_DP1_18_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_18),
  .pullen(`DP1_18_PULLEN),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE)
));
ap_DP1_18_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_18_PINCTRL_0_IE),
  .outen(`DP1_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_18),
  .pad(`DP1_18),
  .default_value(`default_value)));
ap_DP1_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_18_PULLEN),
  .pullsel(`DP1_18_PULLSEL),
  .pad_pullup(`DP1_18)
));
ap_DP1_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_18),
  .pullen(`DP1_18_PULLEN),
  .pullsel(`DP1_18_PULLSEL)
));
ap_DP1_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_18_PULLEN),
  .pullsel(`DP1_18_PULLSEL),
  .pad_pd(`DP1_18)
));
ap_DP1_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_18),
  .pullen(`DP1_18_PULLEN),
  .pullsel(`DP1_18_PULLSEL)
));
ap_DP1_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP1_19),
  .pad_gz(`DP1_19_pad_y)
));
ap_DP1_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP1_19),
  .pad_gz(`DP1_19_pad_y)
));
ap_DP1_19_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_19),
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE)
));
ap_DP1_19_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_19_PINCTRL_0_IE),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_19),
  .pad(`DP1_19),
  .default_value(`default_value)));
ap_DP1_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP1_19),
  .pad_gz(`DP1_19_pad_y)
));
ap_DP1_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_19),
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE)
));
ap_DP1_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_19_PINCTRL_0_IE),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_19),
  .pad(`DP1_19),
  .default_value(`default_value)));
ap_DP1_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_19_OUTFUNC_SEL),
  .gpioouten(`DP1_19_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`DP1_19_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`DP1_19),
  .pad_gz(`DP1_19_pad_y)
));
ap_DP1_19_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_19)
));
ap_DP1_19_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_19),
  .pullen(`DP1_19_PULLEN),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE)
));
ap_DP1_19_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_19_PINCTRL_0_IE),
  .outen(`DP1_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_19),
  .pad(`DP1_19),
  .default_value(`default_value)));
ap_DP1_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_19_PULLEN),
  .pullsel(`DP1_19_PULLSEL),
  .pad_pullup(`DP1_19)
));
ap_DP1_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_19),
  .pullen(`DP1_19_PULLEN),
  .pullsel(`DP1_19_PULLSEL)
));
ap_DP1_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_19_PULLEN),
  .pullsel(`DP1_19_PULLSEL),
  .pad_pd(`DP1_19)
));
ap_DP1_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_19),
  .pullen(`DP1_19_PULLEN),
  .pullsel(`DP1_19_PULLSEL)
));
ap_DP1_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP1_20),
  .pad_gz(`DP1_20_pad_y)
));
ap_DP1_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP1_20),
  .pad_gz(`DP1_20_pad_y)
));
ap_DP1_20_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_20),
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE)
));
ap_DP1_20_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_20_PINCTRL_0_IE),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_20),
  .pad(`DP1_20),
  .default_value(`default_value)));
ap_DP1_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP1_20),
  .pad_gz(`DP1_20_pad_y)
));
ap_DP1_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_20),
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE)
));
ap_DP1_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_20_PINCTRL_0_IE),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_20),
  .pad(`DP1_20),
  .default_value(`default_value)));
ap_DP1_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_20_OUTFUNC_SEL),
  .gpioouten(`DP1_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`DP1_20_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`DP1_20),
  .pad_gz(`DP1_20_pad_y)
));
ap_DP1_20_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_20)
));
ap_DP1_20_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_20),
  .pullen(`DP1_20_PULLEN),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE)
));
ap_DP1_20_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_20_PINCTRL_0_IE),
  .outen(`DP1_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_20),
  .pad(`DP1_20),
  .default_value(`default_value)));
ap_DP1_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_20_PULLEN),
  .pullsel(`DP1_20_PULLSEL),
  .pad_pullup(`DP1_20)
));
ap_DP1_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_20),
  .pullen(`DP1_20_PULLEN),
  .pullsel(`DP1_20_PULLSEL)
));
ap_DP1_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_20_PULLEN),
  .pullsel(`DP1_20_PULLSEL),
  .pad_pd(`DP1_20)
));
ap_DP1_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_20),
  .pullen(`DP1_20_PULLEN),
  .pullsel(`DP1_20_PULLSEL)
));
ap_DP1_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP1_21),
  .pad_gz(`DP1_21_pad_y)
));
ap_DP1_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP1_21),
  .pad_gz(`DP1_21_pad_y)
));
ap_DP1_21_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_21),
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE)
));
ap_DP1_21_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_21_PINCTRL_0_IE),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_21),
  .pad(`DP1_21),
  .default_value(`default_value)));
ap_DP1_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP1_21),
  .pad_gz(`DP1_21_pad_y)
));
ap_DP1_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_21),
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE)
));
ap_DP1_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_21_PINCTRL_0_IE),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_21),
  .pad(`DP1_21),
  .default_value(`default_value)));
ap_DP1_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_21_OUTFUNC_SEL),
  .gpioouten(`DP1_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`DP1_21_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`DP1_21),
  .pad_gz(`DP1_21_pad_y)
));
ap_DP1_21_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_21)
));
ap_DP1_21_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_21),
  .pullen(`DP1_21_PULLEN),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE)
));
ap_DP1_21_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_21_PINCTRL_0_IE),
  .outen(`DP1_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_21),
  .pad(`DP1_21),
  .default_value(`default_value)));
ap_DP1_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_21_PULLEN),
  .pullsel(`DP1_21_PULLSEL),
  .pad_pullup(`DP1_21)
));
ap_DP1_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_21),
  .pullen(`DP1_21_PULLEN),
  .pullsel(`DP1_21_PULLSEL)
));
ap_DP1_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_21_PULLEN),
  .pullsel(`DP1_21_PULLSEL),
  .pad_pd(`DP1_21)
));
ap_DP1_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_21),
  .pullen(`DP1_21_PULLEN),
  .pullsel(`DP1_21_PULLSEL)
));
ap_DP1_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP1_22),
  .pad_gz(`DP1_22_pad_y)
));
ap_DP1_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP1_22),
  .pad_gz(`DP1_22_pad_y)
));
ap_DP1_22_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_22),
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE)
));
ap_DP1_22_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_22_PINCTRL_0_IE),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_22),
  .pad(`DP1_22),
  .default_value(`default_value)));
ap_DP1_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP1_22),
  .pad_gz(`DP1_22_pad_y)
));
ap_DP1_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_22),
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE)
));
ap_DP1_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_22_PINCTRL_0_IE),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_22),
  .pad(`DP1_22),
  .default_value(`default_value)));
ap_DP1_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_22_OUTFUNC_SEL),
  .gpioouten(`DP1_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`DP1_22_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`DP1_22),
  .pad_gz(`DP1_22_pad_y)
));
ap_DP1_22_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_22)
));
ap_DP1_22_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_22),
  .pullen(`DP1_22_PULLEN),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE)
));
ap_DP1_22_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP1_22_PINCTRL_0_IE),
  .outen(`DP1_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_22),
  .pad(`DP1_22),
  .default_value(`default_value)));
ap_DP1_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_22_PULLEN),
  .pullsel(`DP1_22_PULLSEL),
  .pad_pullup(`DP1_22)
));
ap_DP1_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_22),
  .pullen(`DP1_22_PULLEN),
  .pullsel(`DP1_22_PULLSEL)
));
ap_DP1_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_22_PULLEN),
  .pullsel(`DP1_22_PULLSEL),
  .pad_pd(`DP1_22)
));
ap_DP1_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_22),
  .pullen(`DP1_22_PULLEN),
  .pullsel(`DP1_22_PULLSEL)
));
ap_DP1_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP1_23)
));
ap_DP1_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP1_23),
  .pad_gz(`DP1_23_pad_y)
));
ap_DP1_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP1_23)
));
ap_DP1_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP1_23),
  .pad_gz(`DP1_23_pad_y)
));
ap_DP1_23_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_23_PULLEN),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_23)
));
ap_DP1_23_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_23),
  .pullen(`DP1_23_PULLEN),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE)
));
ap_DP1_23_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP1_23_PINCTRL_0_IE),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_23),
  .pad(`DP1_23),
  .default_value(`default_value)));
ap_DP1_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP1_23)
));
ap_DP1_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_23_OUTFUNC_SEL),
  .gpioouten(`DP1_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP1_23_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP1_23),
  .pad_gz(`DP1_23_pad_y)
));
ap_DP1_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_23_PULLEN),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_23)
));
ap_DP1_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_23),
  .pullen(`DP1_23_PULLEN),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE)
));
ap_DP1_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_23_PINCTRL_0_IE),
  .outen(`DP1_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_23),
  .pad(`DP1_23),
  .default_value(`default_value)));
ap_DP1_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_23_PULLEN),
  .pullsel(`DP1_23_PULLSEL),
  .pad_pullup(`DP1_23)
));
ap_DP1_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_23),
  .pullen(`DP1_23_PULLEN),
  .pullsel(`DP1_23_PULLSEL)
));
ap_DP1_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_23_PULLEN),
  .pullsel(`DP1_23_PULLSEL),
  .pad_pd(`DP1_23)
));
ap_DP1_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_23),
  .pullen(`DP1_23_PULLEN),
  .pullsel(`DP1_23_PULLSEL)
));
ap_DP1_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP1_24)
));
ap_DP1_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP1_24),
  .pad_gz(`DP1_24_pad_y)
));
ap_DP1_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP1_24)
));
ap_DP1_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP1_24),
  .pad_gz(`DP1_24_pad_y)
));
ap_DP1_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP1_24)
));
ap_DP1_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL0_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL0_OUT),
  .pad(`DP1_24),
  .pad_gz(`DP1_24_pad_y)
));
ap_DP1_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP1_24)
));
ap_DP1_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_24_OUTFUNC_SEL),
  .gpioouten(`DP1_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP1_24_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP1_24),
  .pad_gz(`DP1_24_pad_y)
));
ap_DP1_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_24_PULLEN),
  .outen(`DP1_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_24)
));
ap_DP1_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_24),
  .pullen(`DP1_24_PULLEN),
  .outen(`DP1_24_GPIO_OUTPUT_ENABLE)
));
ap_DP1_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_24_PINCTRL_0_IE),
  .outen(`DP1_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_24),
  .pad(`DP1_24),
  .default_value(`default_value)));
ap_DP1_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_24_PULLEN),
  .pullsel(`DP1_24_PULLSEL),
  .pad_pullup(`DP1_24)
));
ap_DP1_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_24),
  .pullen(`DP1_24_PULLEN),
  .pullsel(`DP1_24_PULLSEL)
));
ap_DP1_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_24_PULLEN),
  .pullsel(`DP1_24_PULLSEL),
  .pad_pd(`DP1_24)
));
ap_DP1_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_24),
  .pullen(`DP1_24_PULLEN),
  .pullsel(`DP1_24_PULLSEL)
));
ap_DP1_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP1_25)
));
ap_DP1_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP1_25),
  .pad_gz(`DP1_25_pad_y)
));
ap_DP1_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP1_25)
));
ap_DP1_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP1_25),
  .pad_gz(`DP1_25_pad_y)
));
ap_DP1_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP1_25)
));
ap_DP1_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL1_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL1_OUT),
  .pad(`DP1_25),
  .pad_gz(`DP1_25_pad_y)
));
ap_DP1_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP1_25)
));
ap_DP1_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_25_OUTFUNC_SEL),
  .gpioouten(`DP1_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP1_25_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP1_25),
  .pad_gz(`DP1_25_pad_y)
));
ap_DP1_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_25_PULLEN),
  .outen(`DP1_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_25)
));
ap_DP1_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_25),
  .pullen(`DP1_25_PULLEN),
  .outen(`DP1_25_GPIO_OUTPUT_ENABLE)
));
ap_DP1_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_25_PINCTRL_0_IE),
  .outen(`DP1_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_25),
  .pad(`DP1_25),
  .default_value(`default_value)));
ap_DP1_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_25_PULLEN),
  .pullsel(`DP1_25_PULLSEL),
  .pad_pullup(`DP1_25)
));
ap_DP1_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_25),
  .pullen(`DP1_25_PULLEN),
  .pullsel(`DP1_25_PULLSEL)
));
ap_DP1_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_25_PULLEN),
  .pullsel(`DP1_25_PULLSEL),
  .pad_pd(`DP1_25)
));
ap_DP1_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_25),
  .pullen(`DP1_25_PULLEN),
  .pullsel(`DP1_25_PULLSEL)
));
ap_DP1_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP1_26)
));
ap_DP1_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP1_26),
  .pad_gz(`DP1_26_pad_y)
));
ap_DP1_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP1_26)
));
ap_DP1_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP1_26),
  .pad_gz(`DP1_26_pad_y)
));
ap_DP1_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP1_26)
));
ap_DP1_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL2_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL2_OUT),
  .pad(`DP1_26),
  .pad_gz(`DP1_26_pad_y)
));
ap_DP1_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP1_26)
));
ap_DP1_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_26_OUTFUNC_SEL),
  .gpioouten(`DP1_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP1_26_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP1_26),
  .pad_gz(`DP1_26_pad_y)
));
ap_DP1_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_26_PULLEN),
  .outen(`DP1_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_26)
));
ap_DP1_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_26),
  .pullen(`DP1_26_PULLEN),
  .outen(`DP1_26_GPIO_OUTPUT_ENABLE)
));
ap_DP1_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_26_PINCTRL_0_IE),
  .outen(`DP1_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_26),
  .pad(`DP1_26),
  .default_value(`default_value)));
ap_DP1_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_26_PULLEN),
  .pullsel(`DP1_26_PULLSEL),
  .pad_pullup(`DP1_26)
));
ap_DP1_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_26),
  .pullen(`DP1_26_PULLEN),
  .pullsel(`DP1_26_PULLSEL)
));
ap_DP1_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_26_PULLEN),
  .pullsel(`DP1_26_PULLSEL),
  .pad_pd(`DP1_26)
));
ap_DP1_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_26),
  .pullen(`DP1_26_PULLEN),
  .pullsel(`DP1_26_PULLSEL)
));
ap_DP1_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP1_27)
));
ap_DP1_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP1_27),
  .pad_gz(`DP1_27_pad_y)
));
ap_DP1_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP1_27)
));
ap_DP1_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP1_27),
  .pad_gz(`DP1_27_pad_y)
));
ap_DP1_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP1_27)
));
ap_DP1_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`ADC0EXTMUXSEL3_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`ADC0EXTMUXSEL3_OUT),
  .pad(`DP1_27),
  .pad_gz(`DP1_27_pad_y)
));
ap_DP1_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP1_27)
));
ap_DP1_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_27_OUTFUNC_SEL),
  .gpioouten(`DP1_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP1_27_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP1_27),
  .pad_gz(`DP1_27_pad_y)
));
ap_DP1_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_27_PULLEN),
  .outen(`DP1_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_27)
));
ap_DP1_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_27),
  .pullen(`DP1_27_PULLEN),
  .outen(`DP1_27_GPIO_OUTPUT_ENABLE)
));
ap_DP1_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_27_PINCTRL_0_IE),
  .outen(`DP1_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_27),
  .pad(`DP1_27),
  .default_value(`default_value)));
ap_DP1_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_27_PULLEN),
  .pullsel(`DP1_27_PULLSEL),
  .pad_pullup(`DP1_27)
));
ap_DP1_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_27),
  .pullen(`DP1_27_PULLEN),
  .pullsel(`DP1_27_PULLSEL)
));
ap_DP1_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_27_PULLEN),
  .pullsel(`DP1_27_PULLSEL),
  .pad_pd(`DP1_27)
));
ap_DP1_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_27),
  .pullen(`DP1_27_PULLEN),
  .pullsel(`DP1_27_PULLSEL)
));
ap_DP1_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP1_28)
));
ap_DP1_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP1_28),
  .pad_gz(`DP1_28_pad_y)
));
ap_DP1_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP1_28)
));
ap_DP1_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP1_28),
  .pad_gz(`DP1_28_pad_y)
));
ap_DP1_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL0_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL0_OUT),
  .pad(`DP1_28)
));
ap_DP1_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL0_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL0_OUT),
  .pad(`DP1_28),
  .pad_gz(`DP1_28_pad_y)
));
ap_DP1_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP1_28)
));
ap_DP1_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_28_OUTFUNC_SEL),
  .gpioouten(`DP1_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP1_28_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP1_28),
  .pad_gz(`DP1_28_pad_y)
));
ap_DP1_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_28_PULLEN),
  .outen(`DP1_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_28)
));
ap_DP1_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_28),
  .pullen(`DP1_28_PULLEN),
  .outen(`DP1_28_GPIO_OUTPUT_ENABLE)
));
ap_DP1_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_28_PINCTRL_0_IE),
  .outen(`DP1_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_28),
  .pad(`DP1_28),
  .default_value(`default_value)));
ap_DP1_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_28_PULLEN),
  .pullsel(`DP1_28_PULLSEL),
  .pad_pullup(`DP1_28)
));
ap_DP1_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_28),
  .pullen(`DP1_28_PULLEN),
  .pullsel(`DP1_28_PULLSEL)
));
ap_DP1_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_28_PULLEN),
  .pullsel(`DP1_28_PULLSEL),
  .pad_pd(`DP1_28)
));
ap_DP1_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_28),
  .pullen(`DP1_28_PULLEN),
  .pullsel(`DP1_28_PULLSEL)
));
ap_DP1_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP1_29)
));
ap_DP1_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP1_29),
  .pad_gz(`DP1_29_pad_y)
));
ap_DP1_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP1_29)
));
ap_DP1_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP1_29),
  .pad_gz(`DP1_29_pad_y)
));
ap_DP1_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL1_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL1_OUT),
  .pad(`DP1_29)
));
ap_DP1_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL1_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL1_OUT),
  .pad(`DP1_29),
  .pad_gz(`DP1_29_pad_y)
));
ap_DP1_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP1_29)
));
ap_DP1_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_29_OUTFUNC_SEL),
  .gpioouten(`DP1_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP1_29_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP1_29),
  .pad_gz(`DP1_29_pad_y)
));
ap_DP1_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_29_PULLEN),
  .outen(`DP1_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_29)
));
ap_DP1_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_29),
  .pullen(`DP1_29_PULLEN),
  .outen(`DP1_29_GPIO_OUTPUT_ENABLE)
));
ap_DP1_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_29_PINCTRL_0_IE),
  .outen(`DP1_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_29),
  .pad(`DP1_29),
  .default_value(`default_value)));
ap_DP1_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_29_PULLEN),
  .pullsel(`DP1_29_PULLSEL),
  .pad_pullup(`DP1_29)
));
ap_DP1_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_29),
  .pullen(`DP1_29_PULLEN),
  .pullsel(`DP1_29_PULLSEL)
));
ap_DP1_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_29_PULLEN),
  .pullsel(`DP1_29_PULLSEL),
  .pad_pd(`DP1_29)
));
ap_DP1_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_29),
  .pullen(`DP1_29_PULLEN),
  .pullsel(`DP1_29_PULLSEL)
));
ap_DP1_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP1_30)
));
ap_DP1_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP1_30),
  .pad_gz(`DP1_30_pad_y)
));
ap_DP1_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP1_30)
));
ap_DP1_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR14_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR14_OUT),
  .pad(`DP1_30),
  .pad_gz(`DP1_30_pad_y)
));
ap_DP1_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL2_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL2_OUT),
  .pad(`DP1_30)
));
ap_DP1_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL2_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL2_OUT),
  .pad(`DP1_30),
  .pad_gz(`DP1_30_pad_y)
));
ap_DP1_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP1_30)
));
ap_DP1_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_30_OUTFUNC_SEL),
  .gpioouten(`DP1_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP1_30_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP1_30),
  .pad_gz(`DP1_30_pad_y)
));
ap_DP1_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_30_PULLEN),
  .outen(`DP1_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_30)
));
ap_DP1_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_30),
  .pullen(`DP1_30_PULLEN),
  .outen(`DP1_30_GPIO_OUTPUT_ENABLE)
));
ap_DP1_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_30_PINCTRL_0_IE),
  .outen(`DP1_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_30),
  .pad(`DP1_30),
  .default_value(`default_value)));
ap_DP1_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_30_PULLEN),
  .pullsel(`DP1_30_PULLSEL),
  .pad_pullup(`DP1_30)
));
ap_DP1_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_30),
  .pullen(`DP1_30_PULLEN),
  .pullsel(`DP1_30_PULLSEL)
));
ap_DP1_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_30_PULLEN),
  .pullsel(`DP1_30_PULLSEL),
  .pad_pd(`DP1_30)
));
ap_DP1_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_30),
  .pullen(`DP1_30_PULLEN),
  .pullsel(`DP1_30_PULLSEL)
));
ap_DP1_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP1_31)
));
ap_DP1_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP1_31),
  .pad_gz(`DP1_31_pad_y)
));
ap_DP1_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP1_31)
));
ap_DP1_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR15_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR15_OUT),
  .pad(`DP1_31),
  .pad_gz(`DP1_31_pad_y)
));
ap_DP1_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL3_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL3_OUT),
  .pad(`DP1_31)
));
ap_DP1_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL3_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL3_OUT),
  .pad(`DP1_31),
  .pad_gz(`DP1_31_pad_y)
));
ap_DP1_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP1_31)
));
ap_DP1_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP1_31_OUTFUNC_SEL),
  .gpioouten(`DP1_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP1_31_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP1_31),
  .pad_gz(`DP1_31_pad_y)
));
ap_DP1_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP1_31_PULLEN),
  .outen(`DP1_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP1_31)
));
ap_DP1_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP1_31),
  .pullen(`DP1_31_PULLEN),
  .outen(`DP1_31_GPIO_OUTPUT_ENABLE)
));
ap_DP1_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP1_31_PINCTRL_0_IE),
  .outen(`DP1_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP1_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP1_31),
  .pad(`DP1_31),
  .default_value(`default_value)));
ap_DP1_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP1_31_PULLEN),
  .pullsel(`DP1_31_PULLSEL),
  .pad_pullup(`DP1_31)
));
ap_DP1_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP1_31),
  .pullen(`DP1_31_PULLEN),
  .pullsel(`DP1_31_PULLSEL)
));
ap_DP1_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP1_31_PULLEN),
  .pullsel(`DP1_31_PULLSEL),
  .pad_pd(`DP1_31)
));
ap_DP1_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP1_31),
  .pullen(`DP1_31_PULLEN),
  .pullsel(`DP1_31_PULLSEL)
));
ap_DP2_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP2_0)
));
ap_DP2_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP2_0),
  .pad_gz(`DP2_0_pad_y)
));
ap_DP2_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP2_0)
));
ap_DP2_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP2_0),
  .pad_gz(`DP2_0_pad_y)
));
ap_DP2_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP2_0)
));
ap_DP2_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL0_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL0_OUT),
  .pad(`DP2_0),
  .pad_gz(`DP2_0_pad_y)
));
ap_DP2_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP2_0)
));
ap_DP2_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_0_OUTFUNC_SEL),
  .gpioouten(`DP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP2_0_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP2_0),
  .pad_gz(`DP2_0_pad_y)
));
ap_DP2_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_0_PULLEN),
  .outen(`DP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_0)
));
ap_DP2_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_0),
  .pullen(`DP2_0_PULLEN),
  .outen(`DP2_0_GPIO_OUTPUT_ENABLE)
));
ap_DP2_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_0_PINCTRL_0_IE),
  .outen(`DP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_0),
  .pad(`DP2_0),
  .default_value(`default_value)));
ap_DP2_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_0_PULLEN),
  .pullsel(`DP2_0_PULLSEL),
  .pad_pullup(`DP2_0)
));
ap_DP2_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_0),
  .pullen(`DP2_0_PULLEN),
  .pullsel(`DP2_0_PULLSEL)
));
ap_DP2_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_0_PULLEN),
  .pullsel(`DP2_0_PULLSEL),
  .pad_pd(`DP2_0)
));
ap_DP2_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_0),
  .pullen(`DP2_0_PULLEN),
  .pullsel(`DP2_0_PULLSEL)
));
ap_DP2_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP2_1)
));
ap_DP2_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP2_1),
  .pad_gz(`DP2_1_pad_y)
));
ap_DP2_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP2_1)
));
ap_DP2_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP2_1),
  .pad_gz(`DP2_1_pad_y)
));
ap_DP2_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP2_1)
));
ap_DP2_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL1_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL1_OUT),
  .pad(`DP2_1),
  .pad_gz(`DP2_1_pad_y)
));
ap_DP2_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP2_1)
));
ap_DP2_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_1_OUTFUNC_SEL),
  .gpioouten(`DP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP2_1_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP2_1),
  .pad_gz(`DP2_1_pad_y)
));
ap_DP2_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_1_PULLEN),
  .outen(`DP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_1)
));
ap_DP2_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_1),
  .pullen(`DP2_1_PULLEN),
  .outen(`DP2_1_GPIO_OUTPUT_ENABLE)
));
ap_DP2_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_1_PINCTRL_0_IE),
  .outen(`DP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_1),
  .pad(`DP2_1),
  .default_value(`default_value)));
ap_DP2_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_1_PULLEN),
  .pullsel(`DP2_1_PULLSEL),
  .pad_pullup(`DP2_1)
));
ap_DP2_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_1),
  .pullen(`DP2_1_PULLEN),
  .pullsel(`DP2_1_PULLSEL)
));
ap_DP2_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_1_PULLEN),
  .pullsel(`DP2_1_PULLSEL),
  .pad_pd(`DP2_1)
));
ap_DP2_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_1),
  .pullen(`DP2_1_PULLEN),
  .pullsel(`DP2_1_PULLSEL)
));
ap_DP2_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP2_2)
));
ap_DP2_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP2_2),
  .pad_gz(`DP2_2_pad_y)
));
ap_DP2_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP2_2)
));
ap_DP2_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP2_2),
  .pad_gz(`DP2_2_pad_y)
));
ap_DP2_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP2_2)
));
ap_DP2_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL2_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL2_OUT),
  .pad(`DP2_2),
  .pad_gz(`DP2_2_pad_y)
));
ap_DP2_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP2_2)
));
ap_DP2_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_2_OUTFUNC_SEL),
  .gpioouten(`DP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP2_2_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP2_2),
  .pad_gz(`DP2_2_pad_y)
));
ap_DP2_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_2_PULLEN),
  .outen(`DP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_2)
));
ap_DP2_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_2),
  .pullen(`DP2_2_PULLEN),
  .outen(`DP2_2_GPIO_OUTPUT_ENABLE)
));
ap_DP2_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_2_PINCTRL_0_IE),
  .outen(`DP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_2),
  .pad(`DP2_2),
  .default_value(`default_value)));
ap_DP2_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_2_PULLEN),
  .pullsel(`DP2_2_PULLSEL),
  .pad_pullup(`DP2_2)
));
ap_DP2_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_2),
  .pullen(`DP2_2_PULLEN),
  .pullsel(`DP2_2_PULLSEL)
));
ap_DP2_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_2_PULLEN),
  .pullsel(`DP2_2_PULLSEL),
  .pad_pd(`DP2_2)
));
ap_DP2_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_2),
  .pullen(`DP2_2_PULLEN),
  .pullsel(`DP2_2_PULLSEL)
));
ap_DP2_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP2_3)
));
ap_DP2_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP2_3),
  .pad_gz(`DP2_3_pad_y)
));
ap_DP2_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP2_3)
));
ap_DP2_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP2_3),
  .pad_gz(`DP2_3_pad_y)
));
ap_DP2_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP2_3)
));
ap_DP2_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP2_3),
  .pad_gz(`DP2_3_pad_y)
));
ap_DP2_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP2_3)
));
ap_DP2_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_3_OUTFUNC_SEL),
  .gpioouten(`DP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP2_3_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP2_3),
  .pad_gz(`DP2_3_pad_y)
));
ap_DP2_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_3_PULLEN),
  .outen(`DP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_3)
));
ap_DP2_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_3),
  .pullen(`DP2_3_PULLEN),
  .outen(`DP2_3_GPIO_OUTPUT_ENABLE)
));
ap_DP2_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_3_PINCTRL_0_IE),
  .outen(`DP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_3),
  .pad(`DP2_3),
  .default_value(`default_value)));
ap_DP2_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_3_PULLEN),
  .pullsel(`DP2_3_PULLSEL),
  .pad_pullup(`DP2_3)
));
ap_DP2_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_3),
  .pullen(`DP2_3_PULLEN),
  .pullsel(`DP2_3_PULLSEL)
));
ap_DP2_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_3_PULLEN),
  .pullsel(`DP2_3_PULLSEL),
  .pad_pd(`DP2_3)
));
ap_DP2_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_3),
  .pullen(`DP2_3_PULLEN),
  .pullsel(`DP2_3_PULLSEL)
));
ap_DP2_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP2_4)
));
ap_DP2_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP2_4),
  .pad_gz(`DP2_4_pad_y)
));
ap_DP2_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP2_4)
));
ap_DP2_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP2_4),
  .pad_gz(`DP2_4_pad_y)
));
ap_DP2_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP2_4)
));
ap_DP2_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP2_4),
  .pad_gz(`DP2_4_pad_y)
));
ap_DP2_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP2_4)
));
ap_DP2_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_4_OUTFUNC_SEL),
  .gpioouten(`DP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP2_4_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP2_4),
  .pad_gz(`DP2_4_pad_y)
));
ap_DP2_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_4_PULLEN),
  .outen(`DP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_4)
));
ap_DP2_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_4),
  .pullen(`DP2_4_PULLEN),
  .outen(`DP2_4_GPIO_OUTPUT_ENABLE)
));
ap_DP2_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_4_PINCTRL_0_IE),
  .outen(`DP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_4),
  .pad(`DP2_4),
  .default_value(`default_value)));
ap_DP2_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_4_PULLEN),
  .pullsel(`DP2_4_PULLSEL),
  .pad_pullup(`DP2_4)
));
ap_DP2_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_4),
  .pullen(`DP2_4_PULLEN),
  .pullsel(`DP2_4_PULLSEL)
));
ap_DP2_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_4_PULLEN),
  .pullsel(`DP2_4_PULLSEL),
  .pad_pd(`DP2_4)
));
ap_DP2_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_4),
  .pullen(`DP2_4_PULLEN),
  .pullsel(`DP2_4_PULLSEL)
));
ap_DP2_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP2_5)
));
ap_DP2_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP2_5),
  .pad_gz(`DP2_5_pad_y)
));
ap_DP2_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP2_5)
));
ap_DP2_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP2_5),
  .pad_gz(`DP2_5_pad_y)
));
ap_DP2_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP2_5)
));
ap_DP2_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP2_5),
  .pad_gz(`DP2_5_pad_y)
));
ap_DP2_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP2_5)
));
ap_DP2_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_5_OUTFUNC_SEL),
  .gpioouten(`DP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP2_5_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP2_5),
  .pad_gz(`DP2_5_pad_y)
));
ap_DP2_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_5_PULLEN),
  .outen(`DP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_5)
));
ap_DP2_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_5),
  .pullen(`DP2_5_PULLEN),
  .outen(`DP2_5_GPIO_OUTPUT_ENABLE)
));
ap_DP2_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_5_PINCTRL_0_IE),
  .outen(`DP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_5),
  .pad(`DP2_5),
  .default_value(`default_value)));
ap_DP2_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_5_PULLEN),
  .pullsel(`DP2_5_PULLSEL),
  .pad_pullup(`DP2_5)
));
ap_DP2_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_5),
  .pullen(`DP2_5_PULLEN),
  .pullsel(`DP2_5_PULLSEL)
));
ap_DP2_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_5_PULLEN),
  .pullsel(`DP2_5_PULLSEL),
  .pad_pd(`DP2_5)
));
ap_DP2_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_5),
  .pullen(`DP2_5_PULLEN),
  .pullsel(`DP2_5_PULLSEL)
));
ap_DP2_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP2_6)
));
ap_DP2_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP2_6),
  .pad_gz(`DP2_6_pad_y)
));
ap_DP2_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP2_6)
));
ap_DP2_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP2_6),
  .pad_gz(`DP2_6_pad_y)
));
ap_DP2_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP2_6)
));
ap_DP2_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP2_6),
  .pad_gz(`DP2_6_pad_y)
));
ap_DP2_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP2_6)
));
ap_DP2_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_6_OUTFUNC_SEL),
  .gpioouten(`DP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP2_6_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP2_6),
  .pad_gz(`DP2_6_pad_y)
));
ap_DP2_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_6_PULLEN),
  .outen(`DP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_6)
));
ap_DP2_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_6),
  .pullen(`DP2_6_PULLEN),
  .outen(`DP2_6_GPIO_OUTPUT_ENABLE)
));
ap_DP2_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_6_PINCTRL_0_IE),
  .outen(`DP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_6),
  .pad(`DP2_6),
  .default_value(`default_value)));
ap_DP2_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_6_PULLEN),
  .pullsel(`DP2_6_PULLSEL),
  .pad_pullup(`DP2_6)
));
ap_DP2_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_6),
  .pullen(`DP2_6_PULLEN),
  .pullsel(`DP2_6_PULLSEL)
));
ap_DP2_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_6_PULLEN),
  .pullsel(`DP2_6_PULLSEL),
  .pad_pd(`DP2_6)
));
ap_DP2_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_6),
  .pullen(`DP2_6_PULLEN),
  .pullsel(`DP2_6_PULLSEL)
));
ap_DP2_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP2_7)
));
ap_DP2_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP2_7),
  .pad_gz(`DP2_7_pad_y)
));
ap_DP2_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP2_7)
));
ap_DP2_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP2_7),
  .pad_gz(`DP2_7_pad_y)
));
ap_DP2_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP2_7)
));
ap_DP2_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP2_7),
  .pad_gz(`DP2_7_pad_y)
));
ap_DP2_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP2_7)
));
ap_DP2_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_7_OUTFUNC_SEL),
  .gpioouten(`DP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP2_7_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP2_7),
  .pad_gz(`DP2_7_pad_y)
));
ap_DP2_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_7_PULLEN),
  .outen(`DP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_7)
));
ap_DP2_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_7),
  .pullen(`DP2_7_PULLEN),
  .outen(`DP2_7_GPIO_OUTPUT_ENABLE)
));
ap_DP2_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_7_PINCTRL_0_IE),
  .outen(`DP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_7),
  .pad(`DP2_7),
  .default_value(`default_value)));
ap_DP2_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_7_PULLEN),
  .pullsel(`DP2_7_PULLSEL),
  .pad_pullup(`DP2_7)
));
ap_DP2_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_7),
  .pullen(`DP2_7_PULLEN),
  .pullsel(`DP2_7_PULLSEL)
));
ap_DP2_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_7_PULLEN),
  .pullsel(`DP2_7_PULLSEL),
  .pad_pd(`DP2_7)
));
ap_DP2_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_7),
  .pullen(`DP2_7_PULLEN),
  .pullsel(`DP2_7_PULLSEL)
));
ap_DP2_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP2_8)
));
ap_DP2_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP2_8),
  .pad_gz(`DP2_8_pad_y)
));
ap_DP2_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP2_8)
));
ap_DP2_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP2_8),
  .pad_gz(`DP2_8_pad_y)
));
ap_DP2_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP2_8)
));
ap_DP2_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP2_8),
  .pad_gz(`DP2_8_pad_y)
));
ap_DP2_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP2_8)
));
ap_DP2_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_8_OUTFUNC_SEL),
  .gpioouten(`DP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP2_8_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP2_8),
  .pad_gz(`DP2_8_pad_y)
));
ap_DP2_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_8_PULLEN),
  .outen(`DP2_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_8)
));
ap_DP2_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_8),
  .pullen(`DP2_8_PULLEN),
  .outen(`DP2_8_GPIO_OUTPUT_ENABLE)
));
ap_DP2_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_8_PINCTRL_0_IE),
  .outen(`DP2_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_8),
  .pad(`DP2_8),
  .default_value(`default_value)));
ap_DP2_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_8_PULLEN),
  .pullsel(`DP2_8_PULLSEL),
  .pad_pullup(`DP2_8)
));
ap_DP2_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_8),
  .pullen(`DP2_8_PULLEN),
  .pullsel(`DP2_8_PULLSEL)
));
ap_DP2_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_8_PULLEN),
  .pullsel(`DP2_8_PULLSEL),
  .pad_pd(`DP2_8)
));
ap_DP2_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_8),
  .pullen(`DP2_8_PULLEN),
  .pullsel(`DP2_8_PULLSEL)
));
ap_DP2_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP2_9)
));
ap_DP2_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP2_9),
  .pad_gz(`DP2_9_pad_y)
));
ap_DP2_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP2_9)
));
ap_DP2_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP2_9),
  .pad_gz(`DP2_9_pad_y)
));
ap_DP2_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP2_9)
));
ap_DP2_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP2_9),
  .pad_gz(`DP2_9_pad_y)
));
ap_DP2_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP2_9)
));
ap_DP2_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_9_OUTFUNC_SEL),
  .gpioouten(`DP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP2_9_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP2_9),
  .pad_gz(`DP2_9_pad_y)
));
ap_DP2_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_9_PULLEN),
  .outen(`DP2_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_9)
));
ap_DP2_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_9),
  .pullen(`DP2_9_PULLEN),
  .outen(`DP2_9_GPIO_OUTPUT_ENABLE)
));
ap_DP2_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_9_PINCTRL_0_IE),
  .outen(`DP2_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_9),
  .pad(`DP2_9),
  .default_value(`default_value)));
ap_DP2_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_9_PULLEN),
  .pullsel(`DP2_9_PULLSEL),
  .pad_pullup(`DP2_9)
));
ap_DP2_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_9),
  .pullen(`DP2_9_PULLEN),
  .pullsel(`DP2_9_PULLSEL)
));
ap_DP2_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_9_PULLEN),
  .pullsel(`DP2_9_PULLSEL),
  .pad_pd(`DP2_9)
));
ap_DP2_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_9),
  .pullen(`DP2_9_PULLEN),
  .pullsel(`DP2_9_PULLSEL)
));
ap_DP2_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP2_10)
));
ap_DP2_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP2_10),
  .pad_gz(`DP2_10_pad_y)
));
ap_DP2_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP2_10)
));
ap_DP2_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP2_10),
  .pad_gz(`DP2_10_pad_y)
));
ap_DP2_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP2_10)
));
ap_DP2_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP2_10),
  .pad_gz(`DP2_10_pad_y)
));
ap_DP2_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP2_10)
));
ap_DP2_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_10_OUTFUNC_SEL),
  .gpioouten(`DP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP2_10_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP2_10),
  .pad_gz(`DP2_10_pad_y)
));
ap_DP2_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_10_PULLEN),
  .outen(`DP2_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_10)
));
ap_DP2_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_10),
  .pullen(`DP2_10_PULLEN),
  .outen(`DP2_10_GPIO_OUTPUT_ENABLE)
));
ap_DP2_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_10_PINCTRL_0_IE),
  .outen(`DP2_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_10),
  .pad(`DP2_10),
  .default_value(`default_value)));
ap_DP2_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_10_PULLEN),
  .pullsel(`DP2_10_PULLSEL),
  .pad_pullup(`DP2_10)
));
ap_DP2_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_10),
  .pullen(`DP2_10_PULLEN),
  .pullsel(`DP2_10_PULLSEL)
));
ap_DP2_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_10_PULLEN),
  .pullsel(`DP2_10_PULLSEL),
  .pad_pd(`DP2_10)
));
ap_DP2_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_10),
  .pullen(`DP2_10_PULLEN),
  .pullsel(`DP2_10_PULLSEL)
));
ap_DP2_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP2_11)
));
ap_DP2_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP2_11),
  .pad_gz(`DP2_11_pad_y)
));
ap_DP2_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP2_11)
));
ap_DP2_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP2_11),
  .pad_gz(`DP2_11_pad_y)
));
ap_DP2_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP2_11)
));
ap_DP2_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_11_OUTFUNC_SEL),
  .gpioouten(`DP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP2_11_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP2_11),
  .pad_gz(`DP2_11_pad_y)
));
ap_DP2_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_11_PULLEN),
  .outen(`DP2_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_11)
));
ap_DP2_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_11),
  .pullen(`DP2_11_PULLEN),
  .outen(`DP2_11_GPIO_OUTPUT_ENABLE)
));
ap_DP2_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_11_PINCTRL_0_IE),
  .outen(`DP2_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_11),
  .pad(`DP2_11),
  .default_value(`default_value)));
ap_DP2_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_11_PULLEN),
  .pullsel(`DP2_11_PULLSEL),
  .pad_pullup(`DP2_11)
));
ap_DP2_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_11),
  .pullen(`DP2_11_PULLEN),
  .pullsel(`DP2_11_PULLSEL)
));
ap_DP2_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_11_PULLEN),
  .pullsel(`DP2_11_PULLSEL),
  .pad_pd(`DP2_11)
));
ap_DP2_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_11),
  .pullen(`DP2_11_PULLEN),
  .pullsel(`DP2_11_PULLSEL)
));
ap_DP2_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP2_12),
  .pad_gz(`DP2_12_pad_y)
));
ap_DP2_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP2_12),
  .pad_gz(`DP2_12_pad_y)
));
ap_DP2_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_12),
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE)
));
ap_DP2_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_12_PINCTRL_0_IE),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_12),
  .pad(`DP2_12),
  .default_value(`default_value)));
ap_DP2_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP2_12),
  .pad_gz(`DP2_12_pad_y)
));
ap_DP2_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP2_12),
  .pad_gz(`DP2_12_pad_y)
));
ap_DP2_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_12),
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE)
));
ap_DP2_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_12_PINCTRL_0_IE),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_12),
  .pad(`DP2_12),
  .default_value(`default_value)));
ap_DP2_12_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_12_OUTFUNC_SEL),
  .gpioouten(`DP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP2_12_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP2_12),
  .pad_gz(`DP2_12_pad_y)
));
ap_DP2_12_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_12)
));
ap_DP2_12_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_12),
  .pullen(`DP2_12_PULLEN),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE)
));
ap_DP2_12_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_12_PINCTRL_0_IE),
  .outen(`DP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_12),
  .pad(`DP2_12),
  .default_value(`default_value)));
ap_DP2_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_12_PULLEN),
  .pullsel(`DP2_12_PULLSEL),
  .pad_pullup(`DP2_12)
));
ap_DP2_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_12),
  .pullen(`DP2_12_PULLEN),
  .pullsel(`DP2_12_PULLSEL)
));
ap_DP2_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_12_PULLEN),
  .pullsel(`DP2_12_PULLSEL),
  .pad_pd(`DP2_12)
));
ap_DP2_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_12),
  .pullen(`DP2_12_PULLEN),
  .pullsel(`DP2_12_PULLSEL)
));
ap_DP2_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE)
));
ap_DP2_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_13_PINCTRL_0_IE),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_13),
  .pad(`DP2_13),
  .default_value(`default_value)));
ap_DP2_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE)
));
ap_DP2_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_13_PINCTRL_0_IE),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_13),
  .pad(`DP2_13),
  .default_value(`default_value)));
ap_DP2_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE)
));
ap_DP2_13_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_13_PINCTRL_0_IE),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_13),
  .pad(`DP2_13),
  .default_value(`default_value)));
ap_DP2_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_13_OUTFUNC_SEL),
  .gpioouten(`DP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP2_13_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP2_13),
  .pad_gz(`DP2_13_pad_y)
));
ap_DP2_13_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_13)
));
ap_DP2_13_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE)
));
ap_DP2_13_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_13_PINCTRL_0_IE),
  .outen(`DP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_13),
  .pad(`DP2_13),
  .default_value(`default_value)));
ap_DP2_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_13_PULLEN),
  .pullsel(`DP2_13_PULLSEL),
  .pad_pullup(`DP2_13)
));
ap_DP2_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .pullsel(`DP2_13_PULLSEL)
));
ap_DP2_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_13_PULLEN),
  .pullsel(`DP2_13_PULLSEL),
  .pad_pd(`DP2_13)
));
ap_DP2_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_13),
  .pullen(`DP2_13_PULLEN),
  .pullsel(`DP2_13_PULLSEL)
));
ap_DP2_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE)
));
ap_DP2_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_14_PINCTRL_0_IE),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_14),
  .pad(`DP2_14),
  .default_value(`default_value)));
ap_DP2_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE)
));
ap_DP2_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_14_PINCTRL_0_IE),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_14),
  .pad(`DP2_14),
  .default_value(`default_value)));
ap_DP2_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE)
));
ap_DP2_14_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_14_PINCTRL_0_IE),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_14),
  .pad(`DP2_14),
  .default_value(`default_value)));
ap_DP2_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_14_OUTFUNC_SEL),
  .gpioouten(`DP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP2_14_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP2_14),
  .pad_gz(`DP2_14_pad_y)
));
ap_DP2_14_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_14)
));
ap_DP2_14_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE)
));
ap_DP2_14_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_14_PINCTRL_0_IE),
  .outen(`DP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_14),
  .pad(`DP2_14),
  .default_value(`default_value)));
ap_DP2_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_14_PULLEN),
  .pullsel(`DP2_14_PULLSEL),
  .pad_pullup(`DP2_14)
));
ap_DP2_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .pullsel(`DP2_14_PULLSEL)
));
ap_DP2_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_14_PULLEN),
  .pullsel(`DP2_14_PULLSEL),
  .pad_pd(`DP2_14)
));
ap_DP2_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_14),
  .pullen(`DP2_14_PULLEN),
  .pullsel(`DP2_14_PULLSEL)
));
ap_DP2_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE)
));
ap_DP2_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_15_PINCTRL_0_IE),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_15),
  .pad(`DP2_15),
  .default_value(`default_value)));
ap_DP2_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE)
));
ap_DP2_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_15_PINCTRL_0_IE),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_15),
  .pad(`DP2_15),
  .default_value(`default_value)));
ap_DP2_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE)
));
ap_DP2_15_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_15_PINCTRL_0_IE),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_15),
  .pad(`DP2_15),
  .default_value(`default_value)));
ap_DP2_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_15_OUTFUNC_SEL),
  .gpioouten(`DP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP2_15_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP2_15),
  .pad_gz(`DP2_15_pad_y)
));
ap_DP2_15_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_15)
));
ap_DP2_15_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE)
));
ap_DP2_15_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_15_PINCTRL_0_IE),
  .outen(`DP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_15),
  .pad(`DP2_15),
  .default_value(`default_value)));
ap_DP2_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_15_PULLEN),
  .pullsel(`DP2_15_PULLSEL),
  .pad_pullup(`DP2_15)
));
ap_DP2_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .pullsel(`DP2_15_PULLSEL)
));
ap_DP2_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_15_PULLEN),
  .pullsel(`DP2_15_PULLSEL),
  .pad_pd(`DP2_15)
));
ap_DP2_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_15),
  .pullen(`DP2_15_PULLEN),
  .pullsel(`DP2_15_PULLSEL)
));
ap_DP2_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE)
));
ap_DP2_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_16_PINCTRL_0_IE),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_16),
  .pad(`DP2_16),
  .default_value(`default_value)));
ap_DP2_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE)
));
ap_DP2_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_16_PINCTRL_0_IE),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_16),
  .pad(`DP2_16),
  .default_value(`default_value)));
ap_DP2_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE)
));
ap_DP2_16_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_16_PINCTRL_0_IE),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_16),
  .pad(`DP2_16),
  .default_value(`default_value)));
ap_DP2_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_16_OUTFUNC_SEL),
  .gpioouten(`DP2_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP2_16_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP2_16),
  .pad_gz(`DP2_16_pad_y)
));
ap_DP2_16_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_16)
));
ap_DP2_16_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE)
));
ap_DP2_16_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_16_PINCTRL_0_IE),
  .outen(`DP2_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_16),
  .pad(`DP2_16),
  .default_value(`default_value)));
ap_DP2_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_16_PULLEN),
  .pullsel(`DP2_16_PULLSEL),
  .pad_pullup(`DP2_16)
));
ap_DP2_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .pullsel(`DP2_16_PULLSEL)
));
ap_DP2_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_16_PULLEN),
  .pullsel(`DP2_16_PULLSEL),
  .pad_pd(`DP2_16)
));
ap_DP2_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_16),
  .pullen(`DP2_16_PULLEN),
  .pullsel(`DP2_16_PULLSEL)
));
ap_DP2_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE)
));
ap_DP2_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_17_PINCTRL_0_IE),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_17),
  .pad(`DP2_17),
  .default_value(`default_value)));
ap_DP2_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE)
));
ap_DP2_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_17_PINCTRL_0_IE),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_17),
  .pad(`DP2_17),
  .default_value(`default_value)));
ap_DP2_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE)
));
ap_DP2_17_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_17_PINCTRL_0_IE),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_17),
  .pad(`DP2_17),
  .default_value(`default_value)));
ap_DP2_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_17_OUTFUNC_SEL),
  .gpioouten(`DP2_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP2_17_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP2_17),
  .pad_gz(`DP2_17_pad_y)
));
ap_DP2_17_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_17)
));
ap_DP2_17_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE)
));
ap_DP2_17_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_17_PINCTRL_0_IE),
  .outen(`DP2_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_17),
  .pad(`DP2_17),
  .default_value(`default_value)));
ap_DP2_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_17_PULLEN),
  .pullsel(`DP2_17_PULLSEL),
  .pad_pullup(`DP2_17)
));
ap_DP2_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .pullsel(`DP2_17_PULLSEL)
));
ap_DP2_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_17_PULLEN),
  .pullsel(`DP2_17_PULLSEL),
  .pad_pd(`DP2_17)
));
ap_DP2_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_17),
  .pullen(`DP2_17_PULLEN),
  .pullsel(`DP2_17_PULLSEL)
));
ap_DP2_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE)
));
ap_DP2_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_18_PINCTRL_0_IE),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_18),
  .pad(`DP2_18),
  .default_value(`default_value)));
ap_DP2_18_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE)
));
ap_DP2_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_18_PINCTRL_0_IE),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_18),
  .pad(`DP2_18),
  .default_value(`default_value)));
ap_DP2_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE)
));
ap_DP2_18_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_18_PINCTRL_0_IE),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_18),
  .pad(`DP2_18),
  .default_value(`default_value)));
ap_DP2_18_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_18_OUTFUNC_SEL),
  .gpioouten(`DP2_18_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP2_18_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP2_18),
  .pad_gz(`DP2_18_pad_y)
));
ap_DP2_18_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_18)
));
ap_DP2_18_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE)
));
ap_DP2_18_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_18_PINCTRL_0_IE),
  .outen(`DP2_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_18),
  .pad(`DP2_18),
  .default_value(`default_value)));
ap_DP2_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_18_PULLEN),
  .pullsel(`DP2_18_PULLSEL),
  .pad_pullup(`DP2_18)
));
ap_DP2_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .pullsel(`DP2_18_PULLSEL)
));
ap_DP2_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_18_PULLEN),
  .pullsel(`DP2_18_PULLSEL),
  .pad_pd(`DP2_18)
));
ap_DP2_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_18),
  .pullen(`DP2_18_PULLEN),
  .pullsel(`DP2_18_PULLSEL)
));
ap_DP2_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE)
));
ap_DP2_19_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_19_PINCTRL_0_IE),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_19),
  .pad(`DP2_19),
  .default_value(`default_value)));
ap_DP2_19_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE)
));
ap_DP2_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_19_PINCTRL_0_IE),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_19),
  .pad(`DP2_19),
  .default_value(`default_value)));
ap_DP2_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE)
));
ap_DP2_19_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_19_PINCTRL_0_IE),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_19),
  .pad(`DP2_19),
  .default_value(`default_value)));
ap_DP2_19_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_19_OUTFUNC_SEL),
  .gpioouten(`DP2_19_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP2_19_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP2_19),
  .pad_gz(`DP2_19_pad_y)
));
ap_DP2_19_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_19)
));
ap_DP2_19_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE)
));
ap_DP2_19_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_19_PINCTRL_0_IE),
  .outen(`DP2_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_19),
  .pad(`DP2_19),
  .default_value(`default_value)));
ap_DP2_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_19_PULLEN),
  .pullsel(`DP2_19_PULLSEL),
  .pad_pullup(`DP2_19)
));
ap_DP2_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .pullsel(`DP2_19_PULLSEL)
));
ap_DP2_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_19_PULLEN),
  .pullsel(`DP2_19_PULLSEL),
  .pad_pd(`DP2_19)
));
ap_DP2_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_19),
  .pullen(`DP2_19_PULLEN),
  .pullsel(`DP2_19_PULLSEL)
));
ap_DP2_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE)
));
ap_DP2_20_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_20_PINCTRL_0_IE),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_20),
  .pad(`DP2_20),
  .default_value(`default_value)));
ap_DP2_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE)
));
ap_DP2_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_20_PINCTRL_0_IE),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_20),
  .pad(`DP2_20),
  .default_value(`default_value)));
ap_DP2_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE)
));
ap_DP2_20_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_20_PINCTRL_0_IE),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_20),
  .pad(`DP2_20),
  .default_value(`default_value)));
ap_DP2_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_20_OUTFUNC_SEL),
  .gpioouten(`DP2_20_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP2_20_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP2_20),
  .pad_gz(`DP2_20_pad_y)
));
ap_DP2_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_20)
));
ap_DP2_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE)
));
ap_DP2_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_20_PINCTRL_0_IE),
  .outen(`DP2_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_20),
  .pad(`DP2_20),
  .default_value(`default_value)));
ap_DP2_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_20_PULLEN),
  .pullsel(`DP2_20_PULLSEL),
  .pad_pullup(`DP2_20)
));
ap_DP2_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .pullsel(`DP2_20_PULLSEL)
));
ap_DP2_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_20_PULLEN),
  .pullsel(`DP2_20_PULLSEL),
  .pad_pd(`DP2_20)
));
ap_DP2_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_20),
  .pullen(`DP2_20_PULLEN),
  .pullsel(`DP2_20_PULLSEL)
));
ap_DP2_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE)
));
ap_DP2_21_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_21_PINCTRL_0_IE),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_21),
  .pad(`DP2_21),
  .default_value(`default_value)));
ap_DP2_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE)
));
ap_DP2_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_21_PINCTRL_0_IE),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_21),
  .pad(`DP2_21),
  .default_value(`default_value)));
ap_DP2_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE)
));
ap_DP2_21_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_21_PINCTRL_0_IE),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_21),
  .pad(`DP2_21),
  .default_value(`default_value)));
ap_DP2_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_21_OUTFUNC_SEL),
  .gpioouten(`DP2_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP2_21_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP2_21),
  .pad_gz(`DP2_21_pad_y)
));
ap_DP2_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_21)
));
ap_DP2_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE)
));
ap_DP2_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_21_PINCTRL_0_IE),
  .outen(`DP2_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_21),
  .pad(`DP2_21),
  .default_value(`default_value)));
ap_DP2_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_21_PULLEN),
  .pullsel(`DP2_21_PULLSEL),
  .pad_pullup(`DP2_21)
));
ap_DP2_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .pullsel(`DP2_21_PULLSEL)
));
ap_DP2_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_21_PULLEN),
  .pullsel(`DP2_21_PULLSEL),
  .pad_pd(`DP2_21)
));
ap_DP2_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_21),
  .pullen(`DP2_21_PULLEN),
  .pullsel(`DP2_21_PULLSEL)
));
ap_DP2_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE)
));
ap_DP2_22_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_22_PINCTRL_0_IE),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_22),
  .pad(`DP2_22),
  .default_value(`default_value)));
ap_DP2_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE)
));
ap_DP2_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_22_PINCTRL_0_IE),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_22),
  .pad(`DP2_22),
  .default_value(`default_value)));
ap_DP2_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE)
));
ap_DP2_22_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_22_PINCTRL_0_IE),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_22),
  .pad(`DP2_22),
  .default_value(`default_value)));
ap_DP2_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_22_OUTFUNC_SEL),
  .gpioouten(`DP2_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP2_22_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP2_22),
  .pad_gz(`DP2_22_pad_y)
));
ap_DP2_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_22)
));
ap_DP2_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE)
));
ap_DP2_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_22_PINCTRL_0_IE),
  .outen(`DP2_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_22),
  .pad(`DP2_22),
  .default_value(`default_value)));
ap_DP2_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_22_PULLEN),
  .pullsel(`DP2_22_PULLSEL),
  .pad_pullup(`DP2_22)
));
ap_DP2_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .pullsel(`DP2_22_PULLSEL)
));
ap_DP2_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_22_PULLEN),
  .pullsel(`DP2_22_PULLSEL),
  .pad_pd(`DP2_22)
));
ap_DP2_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_22),
  .pullen(`DP2_22_PULLEN),
  .pullsel(`DP2_22_PULLSEL)
));
ap_DP2_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE)
));
ap_DP2_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_23_PINCTRL_0_IE),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_23),
  .pad(`DP2_23),
  .default_value(`default_value)));
ap_DP2_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE)
));
ap_DP2_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_23_PINCTRL_0_IE),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_23),
  .pad(`DP2_23),
  .default_value(`default_value)));
ap_DP2_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE)
));
ap_DP2_23_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_23_PINCTRL_0_IE),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_23),
  .pad(`DP2_23),
  .default_value(`default_value)));
ap_DP2_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_23_OUTFUNC_SEL),
  .gpioouten(`DP2_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP2_23_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP2_23),
  .pad_gz(`DP2_23_pad_y)
));
ap_DP2_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_23)
));
ap_DP2_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE)
));
ap_DP2_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_23_PINCTRL_0_IE),
  .outen(`DP2_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_23),
  .pad(`DP2_23),
  .default_value(`default_value)));
ap_DP2_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_23_PULLEN),
  .pullsel(`DP2_23_PULLSEL),
  .pad_pullup(`DP2_23)
));
ap_DP2_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .pullsel(`DP2_23_PULLSEL)
));
ap_DP2_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_23_PULLEN),
  .pullsel(`DP2_23_PULLSEL),
  .pad_pd(`DP2_23)
));
ap_DP2_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_23),
  .pullen(`DP2_23_PULLEN),
  .pullsel(`DP2_23_PULLSEL)
));
ap_DP2_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE)
));
ap_DP2_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_24_PINCTRL_0_IE),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_24),
  .pad(`DP2_24),
  .default_value(`default_value)));
ap_DP2_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC0_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`ADCSOC0_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC0_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`ADCSOC0_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE)
));
ap_DP2_24_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_24_PINCTRL_0_IE),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_24),
  .pad(`DP2_24),
  .default_value(`default_value)));
ap_DP2_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE)
));
ap_DP2_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_24_PINCTRL_0_IE),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_24),
  .pad(`DP2_24),
  .default_value(`default_value)));
ap_DP2_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE)
));
ap_DP2_24_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_24_PINCTRL_0_IE),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_24),
  .pad(`DP2_24),
  .default_value(`default_value)));
ap_DP2_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_24_OUTFUNC_SEL),
  .gpioouten(`DP2_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP2_24_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP2_24),
  .pad_gz(`DP2_24_pad_y)
));
ap_DP2_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_24)
));
ap_DP2_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE)
));
ap_DP2_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_24_PINCTRL_0_IE),
  .outen(`DP2_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_24),
  .pad(`DP2_24),
  .default_value(`default_value)));
ap_DP2_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_24_PULLEN),
  .pullsel(`DP2_24_PULLSEL),
  .pad_pullup(`DP2_24)
));
ap_DP2_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .pullsel(`DP2_24_PULLSEL)
));
ap_DP2_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_24_PULLEN),
  .pullsel(`DP2_24_PULLSEL),
  .pad_pd(`DP2_24)
));
ap_DP2_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_24),
  .pullen(`DP2_24_PULLEN),
  .pullsel(`DP2_24_PULLSEL)
));
ap_DP2_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE)
));
ap_DP2_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_25_PINCTRL_0_IE),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_25),
  .pad(`DP2_25),
  .default_value(`default_value)));
ap_DP2_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC1_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`ADCSOC1_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC1_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`ADCSOC1_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE)
));
ap_DP2_25_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_25_PINCTRL_0_IE),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_25),
  .pad(`DP2_25),
  .default_value(`default_value)));
ap_DP2_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE)
));
ap_DP2_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_25_PINCTRL_0_IE),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_25),
  .pad(`DP2_25),
  .default_value(`default_value)));
ap_DP2_25_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE)
));
ap_DP2_25_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_25_PINCTRL_0_IE),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_25),
  .pad(`DP2_25),
  .default_value(`default_value)));
ap_DP2_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_25_OUTFUNC_SEL),
  .gpioouten(`DP2_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP2_25_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP2_25),
  .pad_gz(`DP2_25_pad_y)
));
ap_DP2_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_25)
));
ap_DP2_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE)
));
ap_DP2_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_25_PINCTRL_0_IE),
  .outen(`DP2_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_25),
  .pad(`DP2_25),
  .default_value(`default_value)));
ap_DP2_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_25_PULLEN),
  .pullsel(`DP2_25_PULLSEL),
  .pad_pullup(`DP2_25)
));
ap_DP2_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .pullsel(`DP2_25_PULLSEL)
));
ap_DP2_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_25_PULLEN),
  .pullsel(`DP2_25_PULLSEL),
  .pad_pd(`DP2_25)
));
ap_DP2_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_25),
  .pullen(`DP2_25_PULLEN),
  .pullsel(`DP2_25_PULLSEL)
));
ap_DP2_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE)
));
ap_DP2_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_26_PINCTRL_0_IE),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_26),
  .pad(`DP2_26),
  .default_value(`default_value)));
ap_DP2_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE)
));
ap_DP2_26_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_26_PINCTRL_0_IE),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_26),
  .pad(`DP2_26),
  .default_value(`default_value)));
ap_DP2_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE)
));
ap_DP2_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_26_PINCTRL_0_IE),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_26),
  .pad(`DP2_26),
  .default_value(`default_value)));
ap_DP2_26_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE)
));
ap_DP2_26_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_26_PINCTRL_0_IE),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_26),
  .pad(`DP2_26),
  .default_value(`default_value)));
ap_DP2_26_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_26_OUTFUNC_SEL),
  .gpioouten(`DP2_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP2_26_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP2_26),
  .pad_gz(`DP2_26_pad_y)
));
ap_DP2_26_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_26)
));
ap_DP2_26_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE)
));
ap_DP2_26_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_26_PINCTRL_0_IE),
  .outen(`DP2_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_26),
  .pad(`DP2_26),
  .default_value(`default_value)));
ap_DP2_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_26_PULLEN),
  .pullsel(`DP2_26_PULLSEL),
  .pad_pullup(`DP2_26)
));
ap_DP2_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .pullsel(`DP2_26_PULLSEL)
));
ap_DP2_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_26_PULLEN),
  .pullsel(`DP2_26_PULLSEL),
  .pad_pd(`DP2_26)
));
ap_DP2_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_26),
  .pullen(`DP2_26_PULLEN),
  .pullsel(`DP2_26_PULLSEL)
));
ap_DP2_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE)
));
ap_DP2_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_27_PINCTRL_0_IE),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_27),
  .pad(`DP2_27),
  .default_value(`default_value)));
ap_DP2_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE)
));
ap_DP2_27_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_27_PINCTRL_0_IE),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_27),
  .pad(`DP2_27),
  .default_value(`default_value)));
ap_DP2_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE)
));
ap_DP2_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_27_PINCTRL_0_IE),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_27),
  .pad(`DP2_27),
  .default_value(`default_value)));
ap_DP2_27_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE)
));
ap_DP2_27_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_27_PINCTRL_0_IE),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_27),
  .pad(`DP2_27),
  .default_value(`default_value)));
ap_DP2_27_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_27_OUTFUNC_SEL),
  .gpioouten(`DP2_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP2_27_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP2_27),
  .pad_gz(`DP2_27_pad_y)
));
ap_DP2_27_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_27)
));
ap_DP2_27_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE)
));
ap_DP2_27_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_27_PINCTRL_0_IE),
  .outen(`DP2_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_27),
  .pad(`DP2_27),
  .default_value(`default_value)));
ap_DP2_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_27_PULLEN),
  .pullsel(`DP2_27_PULLSEL),
  .pad_pullup(`DP2_27)
));
ap_DP2_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .pullsel(`DP2_27_PULLSEL)
));
ap_DP2_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_27_PULLEN),
  .pullsel(`DP2_27_PULLSEL),
  .pad_pd(`DP2_27)
));
ap_DP2_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_27),
  .pullen(`DP2_27_PULLEN),
  .pullsel(`DP2_27_PULLSEL)
));
ap_DP2_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE)
));
ap_DP2_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_28_PINCTRL_0_IE),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_28),
  .pad(`DP2_28),
  .default_value(`default_value)));
ap_DP2_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE)
));
ap_DP2_28_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_28_PINCTRL_0_IE),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_28),
  .pad(`DP2_28),
  .default_value(`default_value)));
ap_DP2_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE)
));
ap_DP2_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_28_PINCTRL_0_IE),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_28),
  .pad(`DP2_28),
  .default_value(`default_value)));
ap_DP2_28_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE)
));
ap_DP2_28_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_28_PINCTRL_0_IE),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_28),
  .pad(`DP2_28),
  .default_value(`default_value)));
ap_DP2_28_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_28_OUTFUNC_SEL),
  .gpioouten(`DP2_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP2_28_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP2_28),
  .pad_gz(`DP2_28_pad_y)
));
ap_DP2_28_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_28)
));
ap_DP2_28_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE)
));
ap_DP2_28_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_28_PINCTRL_0_IE),
  .outen(`DP2_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_28),
  .pad(`DP2_28),
  .default_value(`default_value)));
ap_DP2_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_28_PULLEN),
  .pullsel(`DP2_28_PULLSEL),
  .pad_pullup(`DP2_28)
));
ap_DP2_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .pullsel(`DP2_28_PULLSEL)
));
ap_DP2_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_28_PULLEN),
  .pullsel(`DP2_28_PULLSEL),
  .pad_pd(`DP2_28)
));
ap_DP2_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_28),
  .pullen(`DP2_28_PULLEN),
  .pullsel(`DP2_28_PULLSEL)
));
ap_DP2_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP2_29),
  .pad_gz(`DP2_29_pad_y)
));
ap_DP2_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`DP2_29),
  .pad_gz(`DP2_29_pad_y)
));
ap_DP2_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE)
));
ap_DP2_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_29_PINCTRL_0_IE),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_29),
  .pad(`DP2_29),
  .default_value(`default_value)));
ap_DP2_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP2_29),
  .pad_gz(`DP2_29_pad_y)
));
ap_DP2_29_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE)
));
ap_DP2_29_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_29_PINCTRL_0_IE),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_29),
  .pad(`DP2_29),
  .default_value(`default_value)));
ap_DP2_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP2_29),
  .pad_gz(`DP2_29_pad_y)
));
ap_DP2_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE)
));
ap_DP2_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_29_PINCTRL_0_IE),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_29),
  .pad(`DP2_29),
  .default_value(`default_value)));
ap_DP2_29_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE)
));
ap_DP2_29_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_29_PINCTRL_0_IE),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_29),
  .pad(`DP2_29),
  .default_value(`default_value)));
ap_DP2_29_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_29_OUTFUNC_SEL),
  .gpioouten(`DP2_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP2_29_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP2_29),
  .pad_gz(`DP2_29_pad_y)
));
ap_DP2_29_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_29)
));
ap_DP2_29_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE)
));
ap_DP2_29_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_29_PINCTRL_0_IE),
  .outen(`DP2_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_29),
  .pad(`DP2_29),
  .default_value(`default_value)));
ap_DP2_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_29_PULLEN),
  .pullsel(`DP2_29_PULLSEL),
  .pad_pullup(`DP2_29)
));
ap_DP2_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .pullsel(`DP2_29_PULLSEL)
));
ap_DP2_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_29_PULLEN),
  .pullsel(`DP2_29_PULLSEL),
  .pad_pd(`DP2_29)
));
ap_DP2_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_29),
  .pullen(`DP2_29_PULLEN),
  .pullsel(`DP2_29_PULLSEL)
));
ap_DP2_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP2_30),
  .pad_gz(`DP2_30_pad_y)
));
ap_DP2_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`DP2_30),
  .pad_gz(`DP2_30_pad_y)
));
ap_DP2_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE)
));
ap_DP2_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_30_PINCTRL_0_IE),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_30),
  .pad(`DP2_30),
  .default_value(`default_value)));
ap_DP2_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP2_30),
  .pad_gz(`DP2_30_pad_y)
));
ap_DP2_30_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE)
));
ap_DP2_30_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_30_PINCTRL_0_IE),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_30),
  .pad(`DP2_30),
  .default_value(`default_value)));
ap_DP2_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP2_30),
  .pad_gz(`DP2_30_pad_y)
));
ap_DP2_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE)
));
ap_DP2_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_30_PINCTRL_0_IE),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_30),
  .pad(`DP2_30),
  .default_value(`default_value)));
ap_DP2_30_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE)
));
ap_DP2_30_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_30_PINCTRL_0_IE),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_30),
  .pad(`DP2_30),
  .default_value(`default_value)));
ap_DP2_30_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_30_OUTFUNC_SEL),
  .gpioouten(`DP2_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP2_30_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP2_30),
  .pad_gz(`DP2_30_pad_y)
));
ap_DP2_30_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_30)
));
ap_DP2_30_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE)
));
ap_DP2_30_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_30_PINCTRL_0_IE),
  .outen(`DP2_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_30),
  .pad(`DP2_30),
  .default_value(`default_value)));
ap_DP2_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_30_PULLEN),
  .pullsel(`DP2_30_PULLSEL),
  .pad_pullup(`DP2_30)
));
ap_DP2_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .pullsel(`DP2_30_PULLSEL)
));
ap_DP2_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_30_PULLEN),
  .pullsel(`DP2_30_PULLSEL),
  .pad_pd(`DP2_30)
));
ap_DP2_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_30),
  .pullen(`DP2_30_PULLEN),
  .pullsel(`DP2_30_PULLSEL)
));
ap_DP2_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP2_31),
  .pad_gz(`DP2_31_pad_y)
));
ap_DP2_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`DP2_31),
  .pad_gz(`DP2_31_pad_y)
));
ap_DP2_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE)
));
ap_DP2_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP2_31_PINCTRL_0_IE),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_31),
  .pad(`DP2_31),
  .default_value(`default_value)));
ap_DP2_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP2_31),
  .pad_gz(`DP2_31_pad_y)
));
ap_DP2_31_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE)
));
ap_DP2_31_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP2_31_PINCTRL_0_IE),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_31),
  .pad(`DP2_31),
  .default_value(`default_value)));
ap_DP2_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP2_31),
  .pad_gz(`DP2_31_pad_y)
));
ap_DP2_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE)
));
ap_DP2_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP2_31_PINCTRL_0_IE),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_31),
  .pad(`DP2_31),
  .default_value(`default_value)));
ap_DP2_31_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE)
));
ap_DP2_31_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP2_31_PINCTRL_0_IE),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_31),
  .pad(`DP2_31),
  .default_value(`default_value)));
ap_DP2_31_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP2_31_OUTFUNC_SEL),
  .gpioouten(`DP2_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP2_31_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP2_31),
  .pad_gz(`DP2_31_pad_y)
));
ap_DP2_31_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP2_31)
));
ap_DP2_31_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE)
));
ap_DP2_31_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP2_31_PINCTRL_0_IE),
  .outen(`DP2_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP2_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP2_31),
  .pad(`DP2_31),
  .default_value(`default_value)));
ap_DP2_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP2_31_PULLEN),
  .pullsel(`DP2_31_PULLSEL),
  .pad_pullup(`DP2_31)
));
ap_DP2_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .pullsel(`DP2_31_PULLSEL)
));
ap_DP2_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP2_31_PULLEN),
  .pullsel(`DP2_31_PULLSEL),
  .pad_pd(`DP2_31)
));
ap_DP2_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP2_31),
  .pullen(`DP2_31_PULLEN),
  .pullsel(`DP2_31_PULLSEL)
));
ap_DP3_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWMSYNCO_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`EPWMSYNCO_OUT),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWMSYNCO_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`EPWMSYNCO_OUT),
  .pad(`DP3_0),
  .pad_gz(`DP3_0_pad_y)
));
ap_DP3_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`DP3_0),
  .pad_gz(`DP3_0_pad_y)
));
ap_DP3_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE)
));
ap_DP3_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_0_PINCTRL_0_IE),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_0),
  .pad(`DP3_0),
  .default_value(`default_value)));
ap_DP3_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP3_0),
  .pad_gz(`DP3_0_pad_y)
));
ap_DP3_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE)
));
ap_DP3_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP3_0_PINCTRL_0_IE),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_0),
  .pad(`DP3_0),
  .default_value(`default_value)));
ap_DP3_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP3_0),
  .pad_gz(`DP3_0_pad_y)
));
ap_DP3_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE)
));
ap_DP3_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_0_PINCTRL_0_IE),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_0),
  .pad(`DP3_0),
  .default_value(`default_value)));
ap_DP3_0_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE)
));
ap_DP3_0_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_0_PINCTRL_0_IE),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_0),
  .pad(`DP3_0),
  .default_value(`default_value)));
ap_DP3_0_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_0_OUTFUNC_SEL),
  .gpioouten(`DP3_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP3_0_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP3_0),
  .pad_gz(`DP3_0_pad_y)
));
ap_DP3_0_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_0)
));
ap_DP3_0_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE)
));
ap_DP3_0_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_0_PINCTRL_0_IE),
  .outen(`DP3_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_0),
  .pad(`DP3_0),
  .default_value(`default_value)));
ap_DP3_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_0_PULLEN),
  .pullsel(`DP3_0_PULLSEL),
  .pad_pullup(`DP3_0)
));
ap_DP3_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .pullsel(`DP3_0_PULLSEL)
));
ap_DP3_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_0_PULLEN),
  .pullsel(`DP3_0_PULLSEL),
  .pad_pd(`DP3_0)
));
ap_DP3_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_0),
  .pullen(`DP3_0_PULLEN),
  .pullsel(`DP3_0_PULLSEL)
));
ap_DP3_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE)
));
ap_DP3_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_1_PINCTRL_0_IE),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_1),
  .pad(`DP3_1),
  .default_value(`default_value)));
ap_DP3_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE)
));
ap_DP3_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_1_PINCTRL_0_IE),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_1),
  .pad(`DP3_1),
  .default_value(`default_value)));
ap_DP3_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD0_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`FSI3TXD0_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD0_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`FSI3TXD0_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE)
));
ap_DP3_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_1_PINCTRL_0_IE),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_1),
  .pad(`DP3_1),
  .default_value(`default_value)));
ap_DP3_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE)
));
ap_DP3_1_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_1_PINCTRL_0_IE),
  .outen(`DP3_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_1),
  .pad(`DP3_1),
  .default_value(`default_value)));
ap_DP3_1_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP3_1)
));
ap_DP3_1_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_1_OUTFUNC_SEL),
  .gpioouten(`DP3_1_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL0_OE),
  .od(`DP3_1_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL0_OUT),
  .pad(`DP3_1),
  .pad_gz(`DP3_1_pad_y)
));
ap_DP3_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_1_PULLEN),
  .pullsel(`DP3_1_PULLSEL),
  .pad_pullup(`DP3_1)
));
ap_DP3_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .pullsel(`DP3_1_PULLSEL)
));
ap_DP3_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_1_PULLEN),
  .pullsel(`DP3_1_PULLSEL),
  .pad_pd(`DP3_1)
));
ap_DP3_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_1),
  .pullen(`DP3_1_PULLEN),
  .pullsel(`DP3_1_PULLSEL)
));
ap_DP3_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE)
));
ap_DP3_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_2_PINCTRL_0_IE),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_2),
  .pad(`DP3_2),
  .default_value(`default_value)));
ap_DP3_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE)
));
ap_DP3_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_2_PINCTRL_0_IE),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_2),
  .pad(`DP3_2),
  .default_value(`default_value)));
ap_DP3_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD1_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`FSI3TXD1_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD1_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`FSI3TXD1_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE)
));
ap_DP3_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_2_PINCTRL_0_IE),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_2),
  .pad(`DP3_2),
  .default_value(`default_value)));
ap_DP3_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE)
));
ap_DP3_2_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_2_PINCTRL_0_IE),
  .outen(`DP3_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_2),
  .pad(`DP3_2),
  .default_value(`default_value)));
ap_DP3_2_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP3_2)
));
ap_DP3_2_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_2_OUTFUNC_SEL),
  .gpioouten(`DP3_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL1_OE),
  .od(`DP3_2_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL1_OUT),
  .pad(`DP3_2),
  .pad_gz(`DP3_2_pad_y)
));
ap_DP3_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_2_PULLEN),
  .pullsel(`DP3_2_PULLSEL),
  .pad_pullup(`DP3_2)
));
ap_DP3_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .pullsel(`DP3_2_PULLSEL)
));
ap_DP3_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_2_PULLEN),
  .pullsel(`DP3_2_PULLSEL),
  .pad_pd(`DP3_2)
));
ap_DP3_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_2),
  .pullen(`DP3_2_PULLEN),
  .pullsel(`DP3_2_PULLSEL)
));
ap_DP3_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE)
));
ap_DP3_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_3_PINCTRL_0_IE),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_3),
  .pad(`DP3_3),
  .default_value(`default_value)));
ap_DP3_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE)
));
ap_DP3_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_3_PINCTRL_0_IE),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_3),
  .pad(`DP3_3),
  .default_value(`default_value)));
ap_DP3_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE)
));
ap_DP3_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_3_PINCTRL_0_IE),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_3),
  .pad(`DP3_3),
  .default_value(`default_value)));
ap_DP3_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE)
));
ap_DP3_3_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_3_PINCTRL_0_IE),
  .outen(`DP3_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_3),
  .pad(`DP3_3),
  .default_value(`default_value)));
ap_DP3_3_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP3_3)
));
ap_DP3_3_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_3_OUTFUNC_SEL),
  .gpioouten(`DP3_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL2_OE),
  .od(`DP3_3_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL2_OUT),
  .pad(`DP3_3),
  .pad_gz(`DP3_3_pad_y)
));
ap_DP3_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_3_PULLEN),
  .pullsel(`DP3_3_PULLSEL),
  .pad_pullup(`DP3_3)
));
ap_DP3_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .pullsel(`DP3_3_PULLSEL)
));
ap_DP3_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_3_PULLEN),
  .pullsel(`DP3_3_PULLSEL),
  .pad_pd(`DP3_3)
));
ap_DP3_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_3),
  .pullen(`DP3_3_PULLEN),
  .pullsel(`DP3_3_PULLSEL)
));
ap_DP3_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE)
));
ap_DP3_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_4_PINCTRL_0_IE),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_4),
  .pad(`DP3_4),
  .default_value(`default_value)));
ap_DP3_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE)
));
ap_DP3_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_4_PINCTRL_0_IE),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_4),
  .pad(`DP3_4),
  .default_value(`default_value)));
ap_DP3_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE)
));
ap_DP3_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_4_PINCTRL_0_IE),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_4),
  .pad(`DP3_4),
  .default_value(`default_value)));
ap_DP3_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE)
));
ap_DP3_4_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_4_PINCTRL_0_IE),
  .outen(`DP3_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_4),
  .pad(`DP3_4),
  .default_value(`default_value)));
ap_DP3_4_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP3_4)
));
ap_DP3_4_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_4_OUTFUNC_SEL),
  .gpioouten(`DP3_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC3EXTMUXSEL3_OE),
  .od(`DP3_4_PINCTRL_0_OD),
  .func_out(`ADC3EXTMUXSEL3_OUT),
  .pad(`DP3_4),
  .pad_gz(`DP3_4_pad_y)
));
ap_DP3_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_4_PULLEN),
  .pullsel(`DP3_4_PULLSEL),
  .pad_pullup(`DP3_4)
));
ap_DP3_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .pullsel(`DP3_4_PULLSEL)
));
ap_DP3_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_4_PULLEN),
  .pullsel(`DP3_4_PULLSEL),
  .pad_pd(`DP3_4)
));
ap_DP3_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_4),
  .pullen(`DP3_4_PULLEN),
  .pullsel(`DP3_4_PULLSEL)
));
ap_DP3_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP3_5),
  .pad_gz(`DP3_5_pad_y)
));
ap_DP3_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE)
));
ap_DP3_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_5_PINCTRL_0_IE),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_5),
  .pad(`DP3_5),
  .default_value(`default_value)));
ap_DP3_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP3_5),
  .pad_gz(`DP3_5_pad_y)
));
ap_DP3_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE)
));
ap_DP3_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_5_PINCTRL_0_IE),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_5),
  .pad(`DP3_5),
  .default_value(`default_value)));
ap_DP3_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP3_5),
  .pad_gz(`DP3_5_pad_y)
));
ap_DP3_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP3_5),
  .pad_gz(`DP3_5_pad_y)
));
ap_DP3_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE)
));
ap_DP3_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_5_PINCTRL_0_IE),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_5),
  .pad(`DP3_5),
  .default_value(`default_value)));
ap_DP3_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_5_OUTFUNC_SEL),
  .gpioouten(`DP3_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP3_5_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP3_5),
  .pad_gz(`DP3_5_pad_y)
));
ap_DP3_5_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_5)
));
ap_DP3_5_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE)
));
ap_DP3_5_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_5_PINCTRL_0_IE),
  .outen(`DP3_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_5),
  .pad(`DP3_5),
  .default_value(`default_value)));
ap_DP3_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_5_PULLEN),
  .pullsel(`DP3_5_PULLSEL),
  .pad_pullup(`DP3_5)
));
ap_DP3_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .pullsel(`DP3_5_PULLSEL)
));
ap_DP3_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_5_PULLEN),
  .pullsel(`DP3_5_PULLSEL),
  .pad_pd(`DP3_5)
));
ap_DP3_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_5),
  .pullen(`DP3_5_PULLEN),
  .pullsel(`DP3_5_PULLSEL)
));
ap_DP3_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP3_6),
  .pad_gz(`DP3_6_pad_y)
));
ap_DP3_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE)
));
ap_DP3_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_6_PINCTRL_0_IE),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_6),
  .pad(`DP3_6),
  .default_value(`default_value)));
ap_DP3_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`DP3_6),
  .pad_gz(`DP3_6_pad_y)
));
ap_DP3_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE)
));
ap_DP3_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_6_PINCTRL_0_IE),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_6),
  .pad(`DP3_6),
  .default_value(`default_value)));
ap_DP3_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP3_6),
  .pad_gz(`DP3_6_pad_y)
));
ap_DP3_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXCLK_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`FSI4TXCLK_OUT),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXCLK_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`FSI4TXCLK_OUT),
  .pad(`DP3_6),
  .pad_gz(`DP3_6_pad_y)
));
ap_DP3_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE)
));
ap_DP3_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_6_PINCTRL_0_IE),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_6),
  .pad(`DP3_6),
  .default_value(`default_value)));
ap_DP3_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_6_OUTFUNC_SEL),
  .gpioouten(`DP3_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP3_6_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP3_6),
  .pad_gz(`DP3_6_pad_y)
));
ap_DP3_6_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_6)
));
ap_DP3_6_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE)
));
ap_DP3_6_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_6_PINCTRL_0_IE),
  .outen(`DP3_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_6),
  .pad(`DP3_6),
  .default_value(`default_value)));
ap_DP3_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_6_PULLEN),
  .pullsel(`DP3_6_PULLSEL),
  .pad_pullup(`DP3_6)
));
ap_DP3_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .pullsel(`DP3_6_PULLSEL)
));
ap_DP3_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_6_PULLEN),
  .pullsel(`DP3_6_PULLSEL),
  .pad_pd(`DP3_6)
));
ap_DP3_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_6),
  .pullen(`DP3_6_PULLEN),
  .pullsel(`DP3_6_PULLSEL)
));
ap_DP3_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP3_7),
  .pad_gz(`DP3_7_pad_y)
));
ap_DP3_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE)
));
ap_DP3_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_7_PINCTRL_0_IE),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_7),
  .pad(`DP3_7),
  .default_value(`default_value)));
ap_DP3_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE)
));
ap_DP3_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_7_PINCTRL_0_IE),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_7),
  .pad(`DP3_7),
  .default_value(`default_value)));
ap_DP3_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP3_7),
  .pad_gz(`DP3_7_pad_y)
));
ap_DP3_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD0_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`FSI4TXD0_OUT),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD0_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`FSI4TXD0_OUT),
  .pad(`DP3_7),
  .pad_gz(`DP3_7_pad_y)
));
ap_DP3_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE)
));
ap_DP3_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_7_PINCTRL_0_IE),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_7),
  .pad(`DP3_7),
  .default_value(`default_value)));
ap_DP3_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_7_OUTFUNC_SEL),
  .gpioouten(`DP3_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP3_7_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP3_7),
  .pad_gz(`DP3_7_pad_y)
));
ap_DP3_7_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_7)
));
ap_DP3_7_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE)
));
ap_DP3_7_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_7_PINCTRL_0_IE),
  .outen(`DP3_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_7),
  .pad(`DP3_7),
  .default_value(`default_value)));
ap_DP3_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_7_PULLEN),
  .pullsel(`DP3_7_PULLSEL),
  .pad_pullup(`DP3_7)
));
ap_DP3_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .pullsel(`DP3_7_PULLSEL)
));
ap_DP3_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_7_PULLEN),
  .pullsel(`DP3_7_PULLSEL),
  .pad_pd(`DP3_7)
));
ap_DP3_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_7),
  .pullen(`DP3_7_PULLEN),
  .pullsel(`DP3_7_PULLSEL)
));
ap_DP3_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP3_8),
  .pad_gz(`DP3_8_pad_y)
));
ap_DP3_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE)
));
ap_DP3_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_8_PINCTRL_0_IE),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_8),
  .pad(`DP3_8),
  .default_value(`default_value)));
ap_DP3_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP3_8),
  .pad_gz(`DP3_8_pad_y)
));
ap_DP3_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE)
));
ap_DP3_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_8_PINCTRL_0_IE),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_8),
  .pad(`DP3_8),
  .default_value(`default_value)));
ap_DP3_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP3_8),
  .pad_gz(`DP3_8_pad_y)
));
ap_DP3_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD1_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`FSI4TXD1_OUT),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD1_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`FSI4TXD1_OUT),
  .pad(`DP3_8),
  .pad_gz(`DP3_8_pad_y)
));
ap_DP3_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE)
));
ap_DP3_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_8_PINCTRL_0_IE),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_8),
  .pad(`DP3_8),
  .default_value(`default_value)));
ap_DP3_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_8_OUTFUNC_SEL),
  .gpioouten(`DP3_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP3_8_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP3_8),
  .pad_gz(`DP3_8_pad_y)
));
ap_DP3_8_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_8)
));
ap_DP3_8_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE)
));
ap_DP3_8_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_8_PINCTRL_0_IE),
  .outen(`DP3_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_8),
  .pad(`DP3_8),
  .default_value(`default_value)));
ap_DP3_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_8_PULLEN),
  .pullsel(`DP3_8_PULLSEL),
  .pad_pullup(`DP3_8)
));
ap_DP3_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .pullsel(`DP3_8_PULLSEL)
));
ap_DP3_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_8_PULLEN),
  .pullsel(`DP3_8_PULLSEL),
  .pad_pd(`DP3_8)
));
ap_DP3_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_8),
  .pullen(`DP3_8_PULLEN),
  .pullsel(`DP3_8_PULLSEL)
));
ap_DP3_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP3_9),
  .pad_gz(`DP3_9_pad_y)
));
ap_DP3_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE)
));
ap_DP3_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_9_PINCTRL_0_IE),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_9),
  .pad(`DP3_9),
  .default_value(`default_value)));
ap_DP3_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP3_9),
  .pad_gz(`DP3_9_pad_y)
));
ap_DP3_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE)
));
ap_DP3_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_9_PINCTRL_0_IE),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_9),
  .pad(`DP3_9),
  .default_value(`default_value)));
ap_DP3_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP3_9),
  .pad_gz(`DP3_9_pad_y)
));
ap_DP3_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXCLK_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`FSI4RXCLK_OUT),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXCLK_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`FSI4RXCLK_OUT),
  .pad(`DP3_9),
  .pad_gz(`DP3_9_pad_y)
));
ap_DP3_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE)
));
ap_DP3_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_9_PINCTRL_0_IE),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_9),
  .pad(`DP3_9),
  .default_value(`default_value)));
ap_DP3_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_9_OUTFUNC_SEL),
  .gpioouten(`DP3_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP3_9_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP3_9),
  .pad_gz(`DP3_9_pad_y)
));
ap_DP3_9_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_9)
));
ap_DP3_9_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE)
));
ap_DP3_9_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_9_PINCTRL_0_IE),
  .outen(`DP3_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_9),
  .pad(`DP3_9),
  .default_value(`default_value)));
ap_DP3_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_9_PULLEN),
  .pullsel(`DP3_9_PULLSEL),
  .pad_pullup(`DP3_9)
));
ap_DP3_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .pullsel(`DP3_9_PULLSEL)
));
ap_DP3_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_9_PULLEN),
  .pullsel(`DP3_9_PULLSEL),
  .pad_pd(`DP3_9)
));
ap_DP3_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_9),
  .pullen(`DP3_9_PULLEN),
  .pullsel(`DP3_9_PULLSEL)
));
ap_DP3_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE)
));
ap_DP3_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_10_PINCTRL_0_IE),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_10),
  .pad(`DP3_10),
  .default_value(`default_value)));
ap_DP3_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE)
));
ap_DP3_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_10_PINCTRL_0_IE),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_10),
  .pad(`DP3_10),
  .default_value(`default_value)));
ap_DP3_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD0_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`FSI4RXD0_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD0_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`FSI4RXD0_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE)
));
ap_DP3_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_10_PINCTRL_0_IE),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_10),
  .pad(`DP3_10),
  .default_value(`default_value)));
ap_DP3_10_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE)
));
ap_DP3_10_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_10_PINCTRL_0_IE),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_10),
  .pad(`DP3_10),
  .default_value(`default_value)));
ap_DP3_10_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_10_OUTFUNC_SEL),
  .gpioouten(`DP3_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP3_10_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP3_10),
  .pad_gz(`DP3_10_pad_y)
));
ap_DP3_10_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_10)
));
ap_DP3_10_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE)
));
ap_DP3_10_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_10_PINCTRL_0_IE),
  .outen(`DP3_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_10),
  .pad(`DP3_10),
  .default_value(`default_value)));
ap_DP3_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_10_PULLEN),
  .pullsel(`DP3_10_PULLSEL),
  .pad_pullup(`DP3_10)
));
ap_DP3_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .pullsel(`DP3_10_PULLSEL)
));
ap_DP3_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_10_PULLEN),
  .pullsel(`DP3_10_PULLSEL),
  .pad_pd(`DP3_10)
));
ap_DP3_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_10),
  .pullen(`DP3_10_PULLEN),
  .pullsel(`DP3_10_PULLSEL)
));
ap_DP3_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE)
));
ap_DP3_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_11_PINCTRL_0_IE),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_11),
  .pad(`DP3_11),
  .default_value(`default_value)));
ap_DP3_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE)
));
ap_DP3_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_11_PINCTRL_0_IE),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_11),
  .pad(`DP3_11),
  .default_value(`default_value)));
ap_DP3_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD1_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`FSI4RXD1_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD1_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`FSI4RXD1_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE)
));
ap_DP3_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_11_PINCTRL_0_IE),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_11),
  .pad(`DP3_11),
  .default_value(`default_value)));
ap_DP3_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE)
));
ap_DP3_11_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_11_PINCTRL_0_IE),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_11),
  .pad(`DP3_11),
  .default_value(`default_value)));
ap_DP3_11_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_11_OUTFUNC_SEL),
  .gpioouten(`DP3_11_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP3_11_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP3_11),
  .pad_gz(`DP3_11_pad_y)
));
ap_DP3_11_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_11)
));
ap_DP3_11_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE)
));
ap_DP3_11_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_11_PINCTRL_0_IE),
  .outen(`DP3_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_11),
  .pad(`DP3_11),
  .default_value(`default_value)));
ap_DP3_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_11_PULLEN),
  .pullsel(`DP3_11_PULLSEL),
  .pad_pullup(`DP3_11)
));
ap_DP3_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .pullsel(`DP3_11_PULLSEL)
));
ap_DP3_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_11_PULLEN),
  .pullsel(`DP3_11_PULLSEL),
  .pad_pd(`DP3_11)
));
ap_DP3_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_11),
  .pullen(`DP3_11_PULLEN),
  .pullsel(`DP3_11_PULLSEL)
));
ap_DP3_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE)
));
ap_DP3_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_12_PINCTRL_0_IE),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_12),
  .pad(`DP3_12),
  .default_value(`default_value)));
ap_DP3_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE)
));
ap_DP3_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_12_PINCTRL_0_IE),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_12),
  .pad(`DP3_12),
  .default_value(`default_value)));
ap_DP3_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXCLK_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`FSI5TXCLK_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXCLK_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`FSI5TXCLK_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE)
));
ap_DP3_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_12_PINCTRL_0_IE),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_12),
  .pad(`DP3_12),
  .default_value(`default_value)));
ap_DP3_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE)
));
ap_DP3_12_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_12_PINCTRL_0_IE),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_12),
  .pad(`DP3_12),
  .default_value(`default_value)));
ap_DP3_12_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_12_OUTFUNC_SEL),
  .gpioouten(`DP3_12_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP3_12_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP3_12),
  .pad_gz(`DP3_12_pad_y)
));
ap_DP3_12_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_12)
));
ap_DP3_12_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE)
));
ap_DP3_12_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_12_PINCTRL_0_IE),
  .outen(`DP3_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_12),
  .pad(`DP3_12),
  .default_value(`default_value)));
ap_DP3_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_12_PULLEN),
  .pullsel(`DP3_12_PULLSEL),
  .pad_pullup(`DP3_12)
));
ap_DP3_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .pullsel(`DP3_12_PULLSEL)
));
ap_DP3_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_12_PULLEN),
  .pullsel(`DP3_12_PULLSEL),
  .pad_pd(`DP3_12)
));
ap_DP3_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_12),
  .pullen(`DP3_12_PULLEN),
  .pullsel(`DP3_12_PULLSEL)
));
ap_DP3_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE)
));
ap_DP3_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_13_PINCTRL_0_IE),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_13),
  .pad(`DP3_13),
  .default_value(`default_value)));
ap_DP3_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE)
));
ap_DP3_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_13_PINCTRL_0_IE),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_13),
  .pad(`DP3_13),
  .default_value(`default_value)));
ap_DP3_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD0_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`FSI5TXD0_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD0_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`FSI5TXD0_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE)
));
ap_DP3_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_13_PINCTRL_0_IE),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_13),
  .pad(`DP3_13),
  .default_value(`default_value)));
ap_DP3_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE)
));
ap_DP3_13_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_13_PINCTRL_0_IE),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_13),
  .pad(`DP3_13),
  .default_value(`default_value)));
ap_DP3_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_13_OUTFUNC_SEL),
  .gpioouten(`DP3_13_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP3_13_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP3_13),
  .pad_gz(`DP3_13_pad_y)
));
ap_DP3_13_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_13)
));
ap_DP3_13_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE)
));
ap_DP3_13_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_13_PINCTRL_0_IE),
  .outen(`DP3_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_13),
  .pad(`DP3_13),
  .default_value(`default_value)));
ap_DP3_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_13_PULLEN),
  .pullsel(`DP3_13_PULLSEL),
  .pad_pullup(`DP3_13)
));
ap_DP3_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .pullsel(`DP3_13_PULLSEL)
));
ap_DP3_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_13_PULLEN),
  .pullsel(`DP3_13_PULLSEL),
  .pad_pd(`DP3_13)
));
ap_DP3_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_13),
  .pullen(`DP3_13_PULLEN),
  .pullsel(`DP3_13_PULLSEL)
));
ap_DP3_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE)
));
ap_DP3_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_14_PINCTRL_0_IE),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_14),
  .pad(`DP3_14),
  .default_value(`default_value)));
ap_DP3_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC2EXTMUXSEL3_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`ADC2EXTMUXSEL3_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD1_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`FSI5TXD1_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD1_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`FSI5TXD1_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE)
));
ap_DP3_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_14_PINCTRL_0_IE),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_14),
  .pad(`DP3_14),
  .default_value(`default_value)));
ap_DP3_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE)
));
ap_DP3_14_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_14_PINCTRL_0_IE),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_14),
  .pad(`DP3_14),
  .default_value(`default_value)));
ap_DP3_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_14_OUTFUNC_SEL),
  .gpioouten(`DP3_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`DP3_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`DP3_14),
  .pad_gz(`DP3_14_pad_y)
));
ap_DP3_14_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_14)
));
ap_DP3_14_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE)
));
ap_DP3_14_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_14_PINCTRL_0_IE),
  .outen(`DP3_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_14),
  .pad(`DP3_14),
  .default_value(`default_value)));
ap_DP3_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_14_PULLEN),
  .pullsel(`DP3_14_PULLSEL),
  .pad_pullup(`DP3_14)
));
ap_DP3_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .pullsel(`DP3_14_PULLSEL)
));
ap_DP3_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_14_PULLEN),
  .pullsel(`DP3_14_PULLSEL),
  .pad_pd(`DP3_14)
));
ap_DP3_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_14),
  .pullen(`DP3_14_PULLEN),
  .pullsel(`DP3_14_PULLSEL)
));
ap_DP3_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE)
));
ap_DP3_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_15_PINCTRL_0_IE),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_15),
  .pad(`DP3_15),
  .default_value(`default_value)));
ap_DP3_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE)
));
ap_DP3_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_15_PINCTRL_0_IE),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_15),
  .pad(`DP3_15),
  .default_value(`default_value)));
ap_DP3_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXCLK_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`FSI5RXCLK_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXCLK_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`FSI5RXCLK_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE)
));
ap_DP3_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_15_PINCTRL_0_IE),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_15),
  .pad(`DP3_15),
  .default_value(`default_value)));
ap_DP3_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE)
));
ap_DP3_15_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_15_PINCTRL_0_IE),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_15),
  .pad(`DP3_15),
  .default_value(`default_value)));
ap_DP3_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_15_OUTFUNC_SEL),
  .gpioouten(`DP3_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`DP3_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`DP3_15),
  .pad_gz(`DP3_15_pad_y)
));
ap_DP3_15_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_15)
));
ap_DP3_15_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE)
));
ap_DP3_15_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_15_PINCTRL_0_IE),
  .outen(`DP3_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_15),
  .pad(`DP3_15),
  .default_value(`default_value)));
ap_DP3_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_15_PULLEN),
  .pullsel(`DP3_15_PULLSEL),
  .pad_pullup(`DP3_15)
));
ap_DP3_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .pullsel(`DP3_15_PULLSEL)
));
ap_DP3_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_15_PULLEN),
  .pullsel(`DP3_15_PULLSEL),
  .pad_pd(`DP3_15)
));
ap_DP3_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_15),
  .pullen(`DP3_15_PULLEN),
  .pullsel(`DP3_15_PULLSEL)
));
ap_DP3_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE)
));
ap_DP3_16_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_16_PINCTRL_0_IE),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_16),
  .pad(`DP3_16),
  .default_value(`default_value)));
ap_DP3_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE)
));
ap_DP3_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_16_PINCTRL_0_IE),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_16),
  .pad(`DP3_16),
  .default_value(`default_value)));
ap_DP3_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD0_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`FSI5RXD0_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD0_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`FSI5RXD0_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE)
));
ap_DP3_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_16_PINCTRL_0_IE),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_16),
  .pad(`DP3_16),
  .default_value(`default_value)));
ap_DP3_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE)
));
ap_DP3_16_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_16_PINCTRL_0_IE),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_16),
  .pad(`DP3_16),
  .default_value(`default_value)));
ap_DP3_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_16_OUTFUNC_SEL),
  .gpioouten(`DP3_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`DP3_16_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`DP3_16),
  .pad_gz(`DP3_16_pad_y)
));
ap_DP3_16_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_16)
));
ap_DP3_16_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE)
));
ap_DP3_16_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_16_PINCTRL_0_IE),
  .outen(`DP3_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_16),
  .pad(`DP3_16),
  .default_value(`default_value)));
ap_DP3_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_16_PULLEN),
  .pullsel(`DP3_16_PULLSEL),
  .pad_pullup(`DP3_16)
));
ap_DP3_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .pullsel(`DP3_16_PULLSEL)
));
ap_DP3_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_16_PULLEN),
  .pullsel(`DP3_16_PULLSEL),
  .pad_pd(`DP3_16)
));
ap_DP3_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_16),
  .pullen(`DP3_16_PULLEN),
  .pullsel(`DP3_16_PULLSEL)
));
ap_DP3_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE)
));
ap_DP3_17_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_17_PINCTRL_0_IE),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_17),
  .pad(`DP3_17),
  .default_value(`default_value)));
ap_DP3_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE)
));
ap_DP3_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_17_PINCTRL_0_IE),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_17),
  .pad(`DP3_17),
  .default_value(`default_value)));
ap_DP3_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD1_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`FSI5RXD1_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD1_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`FSI5RXD1_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE)
));
ap_DP3_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_17_PINCTRL_0_IE),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_17),
  .pad(`DP3_17),
  .default_value(`default_value)));
ap_DP3_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE)
));
ap_DP3_17_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_17_PINCTRL_0_IE),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_17),
  .pad(`DP3_17),
  .default_value(`default_value)));
ap_DP3_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_17_OUTFUNC_SEL),
  .gpioouten(`DP3_17_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`DP3_17_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`DP3_17),
  .pad_gz(`DP3_17_pad_y)
));
ap_DP3_17_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_17)
));
ap_DP3_17_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE)
));
ap_DP3_17_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_17_PINCTRL_0_IE),
  .outen(`DP3_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_17),
  .pad(`DP3_17),
  .default_value(`default_value)));
ap_DP3_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_17_PULLEN),
  .pullsel(`DP3_17_PULLSEL),
  .pad_pullup(`DP3_17)
));
ap_DP3_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .pullsel(`DP3_17_PULLSEL)
));
ap_DP3_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_17_PULLEN),
  .pullsel(`DP3_17_PULLSEL),
  .pad_pd(`DP3_17)
));
ap_DP3_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_17),
  .pullen(`DP3_17_PULLEN),
  .pullsel(`DP3_17_PULLSEL)
));
ap_DP3_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE)
));
ap_DP3_18_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_18_PINCTRL_0_IE),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_18),
  .pad(`DP3_18),
  .default_value(`default_value)));
ap_DP3_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE)
));
ap_DP3_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_18_PINCTRL_0_IE),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_18),
  .pad(`DP3_18),
  .default_value(`default_value)));
ap_DP3_18_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE)
));
ap_DP3_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_18_PINCTRL_0_IE),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_18),
  .pad(`DP3_18),
  .default_value(`default_value)));
ap_DP3_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE)
));
ap_DP3_18_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_18_PINCTRL_0_IE),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_18),
  .pad(`DP3_18),
  .default_value(`default_value)));
ap_DP3_18_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_18_OUTFUNC_SEL),
  .gpioouten(`DP3_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`DP3_18_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`DP3_18),
  .pad_gz(`DP3_18_pad_y)
));
ap_DP3_18_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_18)
));
ap_DP3_18_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE)
));
ap_DP3_18_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_18_PINCTRL_0_IE),
  .outen(`DP3_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_18),
  .pad(`DP3_18),
  .default_value(`default_value)));
ap_DP3_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_18_PULLEN),
  .pullsel(`DP3_18_PULLSEL),
  .pad_pullup(`DP3_18)
));
ap_DP3_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .pullsel(`DP3_18_PULLSEL)
));
ap_DP3_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_18_PULLEN),
  .pullsel(`DP3_18_PULLSEL),
  .pad_pd(`DP3_18)
));
ap_DP3_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_18),
  .pullen(`DP3_18_PULLEN),
  .pullsel(`DP3_18_PULLSEL)
));
ap_DP3_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE)
));
ap_DP3_19_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_19_PINCTRL_0_IE),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_19),
  .pad(`DP3_19),
  .default_value(`default_value)));
ap_DP3_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL0_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL0_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL0_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL0_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE)
));
ap_DP3_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_19_PINCTRL_0_IE),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_19),
  .pad(`DP3_19),
  .default_value(`default_value)));
ap_DP3_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE)
));
ap_DP3_19_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_19_PINCTRL_0_IE),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_19),
  .pad(`DP3_19),
  .default_value(`default_value)));
ap_DP3_19_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_19_OUTFUNC_SEL),
  .gpioouten(`DP3_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`DP3_19_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`DP3_19),
  .pad_gz(`DP3_19_pad_y)
));
ap_DP3_19_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_19)
));
ap_DP3_19_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE)
));
ap_DP3_19_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_19_PINCTRL_0_IE),
  .outen(`DP3_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_19),
  .pad(`DP3_19),
  .default_value(`default_value)));
ap_DP3_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_19_PULLEN),
  .pullsel(`DP3_19_PULLSEL),
  .pad_pullup(`DP3_19)
));
ap_DP3_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .pullsel(`DP3_19_PULLSEL)
));
ap_DP3_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_19_PULLEN),
  .pullsel(`DP3_19_PULLSEL),
  .pad_pd(`DP3_19)
));
ap_DP3_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_19),
  .pullen(`DP3_19_PULLEN),
  .pullsel(`DP3_19_PULLSEL)
));
ap_DP3_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE)
));
ap_DP3_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_20_PINCTRL_0_IE),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_20),
  .pad(`DP3_20),
  .default_value(`default_value)));
ap_DP3_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL1_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL1_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL1_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL1_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE)
));
ap_DP3_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_20_PINCTRL_0_IE),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_20),
  .pad(`DP3_20),
  .default_value(`default_value)));
ap_DP3_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE)
));
ap_DP3_20_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_20_PINCTRL_0_IE),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_20),
  .pad(`DP3_20),
  .default_value(`default_value)));
ap_DP3_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_20_OUTFUNC_SEL),
  .gpioouten(`DP3_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`DP3_20_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`DP3_20),
  .pad_gz(`DP3_20_pad_y)
));
ap_DP3_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_20)
));
ap_DP3_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE)
));
ap_DP3_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_20_PINCTRL_0_IE),
  .outen(`DP3_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_20),
  .pad(`DP3_20),
  .default_value(`default_value)));
ap_DP3_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_20_PULLEN),
  .pullsel(`DP3_20_PULLSEL),
  .pad_pullup(`DP3_20)
));
ap_DP3_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .pullsel(`DP3_20_PULLSEL)
));
ap_DP3_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_20_PULLEN),
  .pullsel(`DP3_20_PULLSEL),
  .pad_pd(`DP3_20)
));
ap_DP3_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_20),
  .pullen(`DP3_20_PULLEN),
  .pullsel(`DP3_20_PULLSEL)
));
ap_DP3_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE)
));
ap_DP3_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_21_PINCTRL_0_IE),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_21),
  .pad(`DP3_21),
  .default_value(`default_value)));
ap_DP3_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL2_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL2_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL2_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL2_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE)
));
ap_DP3_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_21_PINCTRL_0_IE),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_21),
  .pad(`DP3_21),
  .default_value(`default_value)));
ap_DP3_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE)
));
ap_DP3_21_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP3_21_PINCTRL_0_IE),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_21),
  .pad(`DP3_21),
  .default_value(`default_value)));
ap_DP3_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_21_OUTFUNC_SEL),
  .gpioouten(`DP3_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`DP3_21_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`DP3_21),
  .pad_gz(`DP3_21_pad_y)
));
ap_DP3_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_21)
));
ap_DP3_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE)
));
ap_DP3_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_21_PINCTRL_0_IE),
  .outen(`DP3_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_21),
  .pad(`DP3_21),
  .default_value(`default_value)));
ap_DP3_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_21_PULLEN),
  .pullsel(`DP3_21_PULLSEL),
  .pad_pullup(`DP3_21)
));
ap_DP3_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .pullsel(`DP3_21_PULLSEL)
));
ap_DP3_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_21_PULLEN),
  .pullsel(`DP3_21_PULLSEL),
  .pad_pd(`DP3_21)
));
ap_DP3_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_21),
  .pullen(`DP3_21_PULLEN),
  .pullsel(`DP3_21_PULLSEL)
));
ap_DP3_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_22),
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE)
));
ap_DP3_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_22_PINCTRL_0_IE),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_22),
  .pad(`DP3_22),
  .default_value(`default_value)));
ap_DP3_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL3_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL3_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC1EXTMUXSEL3_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`ADC1EXTMUXSEL3_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_22),
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE)
));
ap_DP3_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_22_PINCTRL_0_IE),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_22),
  .pad(`DP3_22),
  .default_value(`default_value)));
ap_DP3_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_22_OUTFUNC_SEL),
  .gpioouten(`DP3_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP3_22_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP3_22),
  .pad_gz(`DP3_22_pad_y)
));
ap_DP3_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_22)
));
ap_DP3_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_22),
  .pullen(`DP3_22_PULLEN),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE)
));
ap_DP3_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_22_PINCTRL_0_IE),
  .outen(`DP3_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_22),
  .pad(`DP3_22),
  .default_value(`default_value)));
ap_DP3_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_22_PULLEN),
  .pullsel(`DP3_22_PULLSEL),
  .pad_pullup(`DP3_22)
));
ap_DP3_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_22),
  .pullen(`DP3_22_PULLEN),
  .pullsel(`DP3_22_PULLSEL)
));
ap_DP3_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_22_PULLEN),
  .pullsel(`DP3_22_PULLSEL),
  .pad_pd(`DP3_22)
));
ap_DP3_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_22),
  .pullen(`DP3_22_PULLEN),
  .pullsel(`DP3_22_PULLSEL)
));
ap_DP3_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE)
));
ap_DP3_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_23_PINCTRL_0_IE),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_23),
  .pad(`DP3_23),
  .default_value(`default_value)));
ap_DP3_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXCLK_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`FSI5TXCLK_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXCLK_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`FSI5TXCLK_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE)
));
ap_DP3_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_23_PINCTRL_0_IE),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_23),
  .pad(`DP3_23),
  .default_value(`default_value)));
ap_DP3_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE)
));
ap_DP3_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_23_PINCTRL_0_IE),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_23),
  .pad(`DP3_23),
  .default_value(`default_value)));
ap_DP3_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_23_OUTFUNC_SEL),
  .gpioouten(`DP3_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP3_23_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP3_23),
  .pad_gz(`DP3_23_pad_y)
));
ap_DP3_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_23)
));
ap_DP3_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE)
));
ap_DP3_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_23_PINCTRL_0_IE),
  .outen(`DP3_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_23),
  .pad(`DP3_23),
  .default_value(`default_value)));
ap_DP3_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_23_PULLEN),
  .pullsel(`DP3_23_PULLSEL),
  .pad_pullup(`DP3_23)
));
ap_DP3_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .pullsel(`DP3_23_PULLSEL)
));
ap_DP3_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_23_PULLEN),
  .pullsel(`DP3_23_PULLSEL),
  .pad_pd(`DP3_23)
));
ap_DP3_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_23),
  .pullen(`DP3_23_PULLEN),
  .pullsel(`DP3_23_PULLSEL)
));
ap_DP3_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE)
));
ap_DP3_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_24_PINCTRL_0_IE),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_24),
  .pad(`DP3_24),
  .default_value(`default_value)));
ap_DP3_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD0_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`FSI5TXD0_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD0_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`FSI5TXD0_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE)
));
ap_DP3_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_24_PINCTRL_0_IE),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_24),
  .pad(`DP3_24),
  .default_value(`default_value)));
ap_DP3_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE)
));
ap_DP3_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_24_PINCTRL_0_IE),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_24),
  .pad(`DP3_24),
  .default_value(`default_value)));
ap_DP3_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_24_OUTFUNC_SEL),
  .gpioouten(`DP3_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP3_24_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP3_24),
  .pad_gz(`DP3_24_pad_y)
));
ap_DP3_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_24)
));
ap_DP3_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE)
));
ap_DP3_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_24_PINCTRL_0_IE),
  .outen(`DP3_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_24),
  .pad(`DP3_24),
  .default_value(`default_value)));
ap_DP3_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_24_PULLEN),
  .pullsel(`DP3_24_PULLSEL),
  .pad_pullup(`DP3_24)
));
ap_DP3_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .pullsel(`DP3_24_PULLSEL)
));
ap_DP3_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_24_PULLEN),
  .pullsel(`DP3_24_PULLSEL),
  .pad_pd(`DP3_24)
));
ap_DP3_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_24),
  .pullen(`DP3_24_PULLEN),
  .pullsel(`DP3_24_PULLSEL)
));
ap_DP3_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE)
));
ap_DP3_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_25_PINCTRL_0_IE),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_25),
  .pad(`DP3_25),
  .default_value(`default_value)));
ap_DP3_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD1_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`FSI5TXD1_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5TXD1_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`FSI5TXD1_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE)
));
ap_DP3_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_25_PINCTRL_0_IE),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_25),
  .pad(`DP3_25),
  .default_value(`default_value)));
ap_DP3_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE)
));
ap_DP3_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_25_PINCTRL_0_IE),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_25),
  .pad(`DP3_25),
  .default_value(`default_value)));
ap_DP3_25_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_25_OUTFUNC_SEL),
  .gpioouten(`DP3_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP3_25_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP3_25),
  .pad_gz(`DP3_25_pad_y)
));
ap_DP3_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_25)
));
ap_DP3_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE)
));
ap_DP3_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_25_PINCTRL_0_IE),
  .outen(`DP3_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_25),
  .pad(`DP3_25),
  .default_value(`default_value)));
ap_DP3_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_25_PULLEN),
  .pullsel(`DP3_25_PULLSEL),
  .pad_pullup(`DP3_25)
));
ap_DP3_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .pullsel(`DP3_25_PULLSEL)
));
ap_DP3_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_25_PULLEN),
  .pullsel(`DP3_25_PULLSEL),
  .pad_pd(`DP3_25)
));
ap_DP3_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_25),
  .pullen(`DP3_25_PULLEN),
  .pullsel(`DP3_25_PULLSEL)
));
ap_DP3_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE)
));
ap_DP3_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_26_PINCTRL_0_IE),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_26),
  .pad(`DP3_26),
  .default_value(`default_value)));
ap_DP3_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXCLK_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`FSI5RXCLK_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXCLK_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`FSI5RXCLK_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE)
));
ap_DP3_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_26_PINCTRL_0_IE),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_26),
  .pad(`DP3_26),
  .default_value(`default_value)));
ap_DP3_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE)
));
ap_DP3_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_26_PINCTRL_0_IE),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_26),
  .pad(`DP3_26),
  .default_value(`default_value)));
ap_DP3_26_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_26_OUTFUNC_SEL),
  .gpioouten(`DP3_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP3_26_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP3_26),
  .pad_gz(`DP3_26_pad_y)
));
ap_DP3_26_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_26)
));
ap_DP3_26_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE)
));
ap_DP3_26_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_26_PINCTRL_0_IE),
  .outen(`DP3_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_26),
  .pad(`DP3_26),
  .default_value(`default_value)));
ap_DP3_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_26_PULLEN),
  .pullsel(`DP3_26_PULLSEL),
  .pad_pullup(`DP3_26)
));
ap_DP3_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .pullsel(`DP3_26_PULLSEL)
));
ap_DP3_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_26_PULLEN),
  .pullsel(`DP3_26_PULLSEL),
  .pad_pd(`DP3_26)
));
ap_DP3_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_26),
  .pullen(`DP3_26_PULLEN),
  .pullsel(`DP3_26_PULLSEL)
));
ap_DP3_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE)
));
ap_DP3_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_27_PINCTRL_0_IE),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_27),
  .pad(`DP3_27),
  .default_value(`default_value)));
ap_DP3_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD0_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`FSI5RXD0_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD0_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`FSI5RXD0_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE)
));
ap_DP3_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_27_PINCTRL_0_IE),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_27),
  .pad(`DP3_27),
  .default_value(`default_value)));
ap_DP3_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE)
));
ap_DP3_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_27_PINCTRL_0_IE),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_27),
  .pad(`DP3_27),
  .default_value(`default_value)));
ap_DP3_27_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29A_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`EPWM29A_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_27_OUTFUNC_SEL),
  .gpioouten(`DP3_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP3_27_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP3_27),
  .pad_gz(`DP3_27_pad_y)
));
ap_DP3_27_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_27)
));
ap_DP3_27_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE)
));
ap_DP3_27_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_27_PINCTRL_0_IE),
  .outen(`DP3_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_27),
  .pad(`DP3_27),
  .default_value(`default_value)));
ap_DP3_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_27_PULLEN),
  .pullsel(`DP3_27_PULLSEL),
  .pad_pullup(`DP3_27)
));
ap_DP3_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .pullsel(`DP3_27_PULLSEL)
));
ap_DP3_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_27_PULLEN),
  .pullsel(`DP3_27_PULLSEL),
  .pad_pd(`DP3_27)
));
ap_DP3_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_27),
  .pullen(`DP3_27_PULLEN),
  .pullsel(`DP3_27_PULLSEL)
));
ap_DP3_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE)
));
ap_DP3_28_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_28_PINCTRL_0_IE),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_28),
  .pad(`DP3_28),
  .default_value(`default_value)));
ap_DP3_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD1_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`FSI5RXD1_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI5RXD1_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`FSI5RXD1_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE)
));
ap_DP3_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_28_PINCTRL_0_IE),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_28),
  .pad(`DP3_28),
  .default_value(`default_value)));
ap_DP3_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM29B_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`EPWM29B_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE)
));
ap_DP3_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_28_PINCTRL_0_IE),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_28),
  .pad(`DP3_28),
  .default_value(`default_value)));
ap_DP3_28_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28B_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`EPWM28B_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_28_OUTFUNC_SEL),
  .gpioouten(`DP3_28_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP3_28_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP3_28),
  .pad_gz(`DP3_28_pad_y)
));
ap_DP3_28_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_28)
));
ap_DP3_28_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE)
));
ap_DP3_28_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP3_28_PINCTRL_0_IE),
  .outen(`DP3_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_28),
  .pad(`DP3_28),
  .default_value(`default_value)));
ap_DP3_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_28_PULLEN),
  .pullsel(`DP3_28_PULLSEL),
  .pad_pullup(`DP3_28)
));
ap_DP3_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .pullsel(`DP3_28_PULLSEL)
));
ap_DP3_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_28_PULLEN),
  .pullsel(`DP3_28_PULLSEL),
  .pad_pd(`DP3_28)
));
ap_DP3_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_28),
  .pullen(`DP3_28_PULLEN),
  .pullsel(`DP3_28_PULLSEL)
));
ap_DP3_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP3_29),
  .pad_gz(`DP3_29_pad_y)
));
ap_DP3_29_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE)
));
ap_DP3_29_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_29_PINCTRL_0_IE),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_29),
  .pad(`DP3_29),
  .default_value(`default_value)));
ap_DP3_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CLK_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`SPI8CLK_OUT),
  .pad(`DP3_29),
  .pad_gz(`DP3_29_pad_y)
));
ap_DP3_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE)
));
ap_DP3_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_29_PINCTRL_0_IE),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_29),
  .pad(`DP3_29),
  .default_value(`default_value)));
ap_DP3_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`DP3_29),
  .pad_gz(`DP3_29_pad_y)
));
ap_DP3_29_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE)
));
ap_DP3_29_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP3_29_PINCTRL_0_IE),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_29),
  .pad(`DP3_29),
  .default_value(`default_value)));
ap_DP3_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP3_29),
  .pad_gz(`DP3_29_pad_y)
));
ap_DP3_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE)
));
ap_DP3_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_29_PINCTRL_0_IE),
  .outen(`DP3_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_29),
  .pad(`DP3_29),
  .default_value(`default_value)));
ap_DP3_29_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP3_29)
));
ap_DP3_29_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_29_OUTFUNC_SEL),
  .gpioouten(`DP3_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM28A_OE),
  .od(`DP3_29_PINCTRL_0_OD),
  .func_out(`EPWM28A_OUT),
  .pad(`DP3_29),
  .pad_gz(`DP3_29_pad_y)
));
ap_DP3_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_29_PULLEN),
  .pullsel(`DP3_29_PULLSEL),
  .pad_pullup(`DP3_29)
));
ap_DP3_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .pullsel(`DP3_29_PULLSEL)
));
ap_DP3_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_29_PULLEN),
  .pullsel(`DP3_29_PULLSEL),
  .pad_pd(`DP3_29)
));
ap_DP3_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_29),
  .pullen(`DP3_29_PULLEN),
  .pullsel(`DP3_29_PULLSEL)
));
ap_DP3_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP3_30),
  .pad_gz(`DP3_30_pad_y)
));
ap_DP3_30_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE)
));
ap_DP3_30_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_30_PINCTRL_0_IE),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_30),
  .pad(`DP3_30),
  .default_value(`default_value)));
ap_DP3_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8PICO_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`SPI8PICO_OUT),
  .pad(`DP3_30),
  .pad_gz(`DP3_30_pad_y)
));
ap_DP3_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE)
));
ap_DP3_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_30_PINCTRL_0_IE),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_30),
  .pad(`DP3_30),
  .default_value(`default_value)));
ap_DP3_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`DP3_30),
  .pad_gz(`DP3_30_pad_y)
));
ap_DP3_30_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE)
));
ap_DP3_30_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP3_30_PINCTRL_0_IE),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_30),
  .pad(`DP3_30),
  .default_value(`default_value)));
ap_DP3_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP3_30),
  .pad_gz(`DP3_30_pad_y)
));
ap_DP3_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE)
));
ap_DP3_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_30_PINCTRL_0_IE),
  .outen(`DP3_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_30),
  .pad(`DP3_30),
  .default_value(`default_value)));
ap_DP3_30_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP3_30)
));
ap_DP3_30_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_30_OUTFUNC_SEL),
  .gpioouten(`DP3_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27B_OE),
  .od(`DP3_30_PINCTRL_0_OD),
  .func_out(`EPWM27B_OUT),
  .pad(`DP3_30),
  .pad_gz(`DP3_30_pad_y)
));
ap_DP3_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_30_PULLEN),
  .pullsel(`DP3_30_PULLSEL),
  .pad_pullup(`DP3_30)
));
ap_DP3_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .pullsel(`DP3_30_PULLSEL)
));
ap_DP3_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_30_PULLEN),
  .pullsel(`DP3_30_PULLSEL),
  .pad_pd(`DP3_30)
));
ap_DP3_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_30),
  .pullen(`DP3_30_PULLEN),
  .pullsel(`DP3_30_PULLSEL)
));
ap_DP3_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP3_31),
  .pad_gz(`DP3_31_pad_y)
));
ap_DP3_31_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE)
));
ap_DP3_31_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP3_31_PINCTRL_0_IE),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_31),
  .pad(`DP3_31),
  .default_value(`default_value)));
ap_DP3_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8POCI_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`SPI8POCI_OUT),
  .pad(`DP3_31),
  .pad_gz(`DP3_31_pad_y)
));
ap_DP3_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE)
));
ap_DP3_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP3_31_PINCTRL_0_IE),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_31),
  .pad(`DP3_31),
  .default_value(`default_value)));
ap_DP3_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`DP3_31),
  .pad_gz(`DP3_31_pad_y)
));
ap_DP3_31_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE)
));
ap_DP3_31_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP3_31_PINCTRL_0_IE),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_31),
  .pad(`DP3_31),
  .default_value(`default_value)));
ap_DP3_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP3_31),
  .pad_gz(`DP3_31_pad_y)
));
ap_DP3_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE)
));
ap_DP3_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP3_31_PINCTRL_0_IE),
  .outen(`DP3_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP3_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP3_31),
  .pad(`DP3_31),
  .default_value(`default_value)));
ap_DP3_31_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP3_31)
));
ap_DP3_31_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP3_31_OUTFUNC_SEL),
  .gpioouten(`DP3_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM27A_OE),
  .od(`DP3_31_PINCTRL_0_OD),
  .func_out(`EPWM27A_OUT),
  .pad(`DP3_31),
  .pad_gz(`DP3_31_pad_y)
));
ap_DP3_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP3_31_PULLEN),
  .pullsel(`DP3_31_PULLSEL),
  .pad_pullup(`DP3_31)
));
ap_DP3_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .pullsel(`DP3_31_PULLSEL)
));
ap_DP3_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP3_31_PULLEN),
  .pullsel(`DP3_31_PULLSEL),
  .pad_pd(`DP3_31)
));
ap_DP3_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP3_31),
  .pullen(`DP3_31_PULLEN),
  .pullsel(`DP3_31_PULLSEL)
));
ap_DP4_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP4_0),
  .pad_gz(`DP4_0_pad_y)
));
ap_DP4_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE)
));
ap_DP4_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_0_PINCTRL_0_IE),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_0),
  .pad(`DP4_0),
  .default_value(`default_value)));
ap_DP4_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS0_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`SPI8CS0_OUT),
  .pad(`DP4_0),
  .pad_gz(`DP4_0_pad_y)
));
ap_DP4_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE)
));
ap_DP4_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_0_PINCTRL_0_IE),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_0),
  .pad(`DP4_0),
  .default_value(`default_value)));
ap_DP4_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`DP4_0),
  .pad_gz(`DP4_0_pad_y)
));
ap_DP4_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE)
));
ap_DP4_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_0_PINCTRL_0_IE),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_0),
  .pad(`DP4_0),
  .default_value(`default_value)));
ap_DP4_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP4_0),
  .pad_gz(`DP4_0_pad_y)
));
ap_DP4_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE)
));
ap_DP4_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_0_PINCTRL_0_IE),
  .outen(`DP4_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_0),
  .pad(`DP4_0),
  .default_value(`default_value)));
ap_DP4_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP4_0)
));
ap_DP4_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_0_OUTFUNC_SEL),
  .gpioouten(`DP4_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP4_0_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP4_0),
  .pad_gz(`DP4_0_pad_y)
));
ap_DP4_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_0_PULLEN),
  .pullsel(`DP4_0_PULLSEL),
  .pad_pullup(`DP4_0)
));
ap_DP4_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .pullsel(`DP4_0_PULLSEL)
));
ap_DP4_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_0_PULLEN),
  .pullsel(`DP4_0_PULLSEL),
  .pad_pd(`DP4_0)
));
ap_DP4_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_0),
  .pullen(`DP4_0_PULLEN),
  .pullsel(`DP4_0_PULLSEL)
));
ap_DP4_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP4_1),
  .pad_gz(`DP4_1_pad_y)
));
ap_DP4_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE)
));
ap_DP4_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_1_PINCTRL_0_IE),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_1),
  .pad(`DP4_1),
  .default_value(`default_value)));
ap_DP4_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS1_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`SPI8CS1_OUT),
  .pad(`DP4_1),
  .pad_gz(`DP4_1_pad_y)
));
ap_DP4_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE)
));
ap_DP4_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_1_PINCTRL_0_IE),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_1),
  .pad(`DP4_1),
  .default_value(`default_value)));
ap_DP4_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`DP4_1),
  .pad_gz(`DP4_1_pad_y)
));
ap_DP4_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE)
));
ap_DP4_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_1_PINCTRL_0_IE),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_1),
  .pad(`DP4_1),
  .default_value(`default_value)));
ap_DP4_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP4_1),
  .pad_gz(`DP4_1_pad_y)
));
ap_DP4_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE)
));
ap_DP4_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_1_PINCTRL_0_IE),
  .outen(`DP4_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_1),
  .pad(`DP4_1),
  .default_value(`default_value)));
ap_DP4_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP4_1)
));
ap_DP4_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_1_OUTFUNC_SEL),
  .gpioouten(`DP4_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP4_1_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP4_1),
  .pad_gz(`DP4_1_pad_y)
));
ap_DP4_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_1_PULLEN),
  .pullsel(`DP4_1_PULLSEL),
  .pad_pullup(`DP4_1)
));
ap_DP4_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .pullsel(`DP4_1_PULLSEL)
));
ap_DP4_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_1_PULLEN),
  .pullsel(`DP4_1_PULLSEL),
  .pad_pd(`DP4_1)
));
ap_DP4_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_1),
  .pullen(`DP4_1_PULLEN),
  .pullsel(`DP4_1_PULLSEL)
));
ap_DP4_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP4_2),
  .pad_gz(`DP4_2_pad_y)
));
ap_DP4_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE)
));
ap_DP4_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_2_PINCTRL_0_IE),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_2),
  .pad(`DP4_2),
  .default_value(`default_value)));
ap_DP4_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS2_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`SPI8CS2_OUT),
  .pad(`DP4_2),
  .pad_gz(`DP4_2_pad_y)
));
ap_DP4_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE)
));
ap_DP4_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_2_PINCTRL_0_IE),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_2),
  .pad(`DP4_2),
  .default_value(`default_value)));
ap_DP4_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`DP4_2),
  .pad_gz(`DP4_2_pad_y)
));
ap_DP4_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE)
));
ap_DP4_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_2_PINCTRL_0_IE),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_2),
  .pad(`DP4_2),
  .default_value(`default_value)));
ap_DP4_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`DP4_2),
  .pad_gz(`DP4_2_pad_y)
));
ap_DP4_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE)
));
ap_DP4_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_2_PINCTRL_0_IE),
  .outen(`DP4_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_2),
  .pad(`DP4_2),
  .default_value(`default_value)));
ap_DP4_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP4_2)
));
ap_DP4_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_2_OUTFUNC_SEL),
  .gpioouten(`DP4_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP4_2_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP4_2),
  .pad_gz(`DP4_2_pad_y)
));
ap_DP4_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_2_PULLEN),
  .pullsel(`DP4_2_PULLSEL),
  .pad_pullup(`DP4_2)
));
ap_DP4_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .pullsel(`DP4_2_PULLSEL)
));
ap_DP4_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_2_PULLEN),
  .pullsel(`DP4_2_PULLSEL),
  .pad_pd(`DP4_2)
));
ap_DP4_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_2),
  .pullen(`DP4_2_PULLEN),
  .pullsel(`DP4_2_PULLSEL)
));
ap_DP4_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP4_3),
  .pad_gz(`DP4_3_pad_y)
));
ap_DP4_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE)
));
ap_DP4_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_3_PINCTRL_0_IE),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_3),
  .pad(`DP4_3),
  .default_value(`default_value)));
ap_DP4_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS3_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`SPI8CS3_OUT),
  .pad(`DP4_3),
  .pad_gz(`DP4_3_pad_y)
));
ap_DP4_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE)
));
ap_DP4_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_3_PINCTRL_0_IE),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_3),
  .pad(`DP4_3),
  .default_value(`default_value)));
ap_DP4_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`DP4_3),
  .pad_gz(`DP4_3_pad_y)
));
ap_DP4_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE)
));
ap_DP4_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_3_PINCTRL_0_IE),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_3),
  .pad(`DP4_3),
  .default_value(`default_value)));
ap_DP4_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`DP4_3),
  .pad_gz(`DP4_3_pad_y)
));
ap_DP4_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE)
));
ap_DP4_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_3_PINCTRL_0_IE),
  .outen(`DP4_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_3),
  .pad(`DP4_3),
  .default_value(`default_value)));
ap_DP4_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP4_3)
));
ap_DP4_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_3_OUTFUNC_SEL),
  .gpioouten(`DP4_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP4_3_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP4_3),
  .pad_gz(`DP4_3_pad_y)
));
ap_DP4_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_3_PULLEN),
  .pullsel(`DP4_3_PULLSEL),
  .pad_pullup(`DP4_3)
));
ap_DP4_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .pullsel(`DP4_3_PULLSEL)
));
ap_DP4_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_3_PULLEN),
  .pullsel(`DP4_3_PULLSEL),
  .pad_pd(`DP4_3)
));
ap_DP4_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_3),
  .pullen(`DP4_3_PULLEN),
  .pullsel(`DP4_3_PULLSEL)
));
ap_DP4_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP4_4),
  .pad_gz(`DP4_4_pad_y)
));
ap_DP4_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE)
));
ap_DP4_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_4_PINCTRL_0_IE),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_4),
  .pad(`DP4_4),
  .default_value(`default_value)));
ap_DP4_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`DP4_4),
  .pad_gz(`DP4_4_pad_y)
));
ap_DP4_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE)
));
ap_DP4_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_4_PINCTRL_0_IE),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_4),
  .pad(`DP4_4),
  .default_value(`default_value)));
ap_DP4_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`DP4_4),
  .pad_gz(`DP4_4_pad_y)
));
ap_DP4_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE)
));
ap_DP4_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_4_PINCTRL_0_IE),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_4),
  .pad(`DP4_4),
  .default_value(`default_value)));
ap_DP4_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP4_4),
  .pad_gz(`DP4_4_pad_y)
));
ap_DP4_4_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_4_OUTFUNC_SEL),
  .gpioouten(`DP4_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_4_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_4),
  .pad_gz(`DP4_4_pad_y)
));
ap_DP4_4_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_4)
));
ap_DP4_4_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE)
));
ap_DP4_4_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_4_PINCTRL_0_IE),
  .outen(`DP4_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_4),
  .pad(`DP4_4),
  .default_value(`default_value)));
ap_DP4_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_4_PULLEN),
  .pullsel(`DP4_4_PULLSEL),
  .pad_pullup(`DP4_4)
));
ap_DP4_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .pullsel(`DP4_4_PULLSEL)
));
ap_DP4_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_4_PULLEN),
  .pullsel(`DP4_4_PULLSEL),
  .pad_pd(`DP4_4)
));
ap_DP4_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_4),
  .pullen(`DP4_4_PULLEN),
  .pullsel(`DP4_4_PULLSEL)
));
ap_DP4_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP4_5),
  .pad_gz(`DP4_5_pad_y)
));
ap_DP4_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE)
));
ap_DP4_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_5_PINCTRL_0_IE),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_5),
  .pad(`DP4_5),
  .default_value(`default_value)));
ap_DP4_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP4_5),
  .pad_gz(`DP4_5_pad_y)
));
ap_DP4_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE)
));
ap_DP4_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_5_PINCTRL_0_IE),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_5),
  .pad(`DP4_5),
  .default_value(`default_value)));
ap_DP4_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`DP4_5),
  .pad_gz(`DP4_5_pad_y)
));
ap_DP4_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE)
));
ap_DP4_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_5_PINCTRL_0_IE),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_5),
  .pad(`DP4_5),
  .default_value(`default_value)));
ap_DP4_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP4_5),
  .pad_gz(`DP4_5_pad_y)
));
ap_DP4_5_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_5_OUTFUNC_SEL),
  .gpioouten(`DP4_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_5_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_5),
  .pad_gz(`DP4_5_pad_y)
));
ap_DP4_5_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_5)
));
ap_DP4_5_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE)
));
ap_DP4_5_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_5_PINCTRL_0_IE),
  .outen(`DP4_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_5),
  .pad(`DP4_5),
  .default_value(`default_value)));
ap_DP4_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_5_PULLEN),
  .pullsel(`DP4_5_PULLSEL),
  .pad_pullup(`DP4_5)
));
ap_DP4_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .pullsel(`DP4_5_PULLSEL)
));
ap_DP4_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_5_PULLEN),
  .pullsel(`DP4_5_PULLSEL),
  .pad_pd(`DP4_5)
));
ap_DP4_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_5),
  .pullen(`DP4_5_PULLEN),
  .pullsel(`DP4_5_PULLSEL)
));
ap_DP4_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXCLK_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`RGMII1TXCLK_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXCLK_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`RGMII1TXCLK_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE)
));
ap_DP4_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_6_PINCTRL_0_IE),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_6),
  .pad(`DP4_6),
  .default_value(`default_value)));
ap_DP4_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE)
));
ap_DP4_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_6_PINCTRL_0_IE),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_6),
  .pad(`DP4_6),
  .default_value(`default_value)));
ap_DP4_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE)
));
ap_DP4_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_6_PINCTRL_0_IE),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_6),
  .pad(`DP4_6),
  .default_value(`default_value)));
ap_DP4_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE)
));
ap_DP4_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_6_PINCTRL_0_IE),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_6),
  .pad(`DP4_6),
  .default_value(`default_value)));
ap_DP4_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE)
));
ap_DP4_6_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_6_PINCTRL_0_IE),
  .outen(`DP4_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_6),
  .pad(`DP4_6),
  .default_value(`default_value)));
ap_DP4_6_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP4_6)
));
ap_DP4_6_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_6_OUTFUNC_SEL),
  .gpioouten(`DP4_6_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP4_6_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP4_6),
  .pad_gz(`DP4_6_pad_y)
));
ap_DP4_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_6_PULLEN),
  .pullsel(`DP4_6_PULLSEL),
  .pad_pullup(`DP4_6)
));
ap_DP4_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .pullsel(`DP4_6_PULLSEL)
));
ap_DP4_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_6_PULLEN),
  .pullsel(`DP4_6_PULLSEL),
  .pad_pd(`DP4_6)
));
ap_DP4_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_6),
  .pullen(`DP4_6_PULLEN),
  .pullsel(`DP4_6_PULLSEL)
));
ap_DP4_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD0_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`RGMII1TXD0_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD0_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`RGMII1TXD0_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE)
));
ap_DP4_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_7_PINCTRL_0_IE),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_7),
  .pad(`DP4_7),
  .default_value(`default_value)));
ap_DP4_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE)
));
ap_DP4_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_7_PINCTRL_0_IE),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_7),
  .pad(`DP4_7),
  .default_value(`default_value)));
ap_DP4_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE)
));
ap_DP4_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_7_PINCTRL_0_IE),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_7),
  .pad(`DP4_7),
  .default_value(`default_value)));
ap_DP4_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE)
));
ap_DP4_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_7_PINCTRL_0_IE),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_7),
  .pad(`DP4_7),
  .default_value(`default_value)));
ap_DP4_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE)
));
ap_DP4_7_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_7_PINCTRL_0_IE),
  .outen(`DP4_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_7),
  .pad(`DP4_7),
  .default_value(`default_value)));
ap_DP4_7_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP4_7)
));
ap_DP4_7_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_7_OUTFUNC_SEL),
  .gpioouten(`DP4_7_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP4_7_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP4_7),
  .pad_gz(`DP4_7_pad_y)
));
ap_DP4_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_7_PULLEN),
  .pullsel(`DP4_7_PULLSEL),
  .pad_pullup(`DP4_7)
));
ap_DP4_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .pullsel(`DP4_7_PULLSEL)
));
ap_DP4_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_7_PULLEN),
  .pullsel(`DP4_7_PULLSEL),
  .pad_pd(`DP4_7)
));
ap_DP4_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_7),
  .pullen(`DP4_7_PULLEN),
  .pullsel(`DP4_7_PULLSEL)
));
ap_DP4_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD1_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`RGMII1TXD1_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD1_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`RGMII1TXD1_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE)
));
ap_DP4_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_8_PINCTRL_0_IE),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_8),
  .pad(`DP4_8),
  .default_value(`default_value)));
ap_DP4_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE)
));
ap_DP4_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_8_PINCTRL_0_IE),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_8),
  .pad(`DP4_8),
  .default_value(`default_value)));
ap_DP4_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE)
));
ap_DP4_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_8_PINCTRL_0_IE),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_8),
  .pad(`DP4_8),
  .default_value(`default_value)));
ap_DP4_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE)
));
ap_DP4_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_8_PINCTRL_0_IE),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_8),
  .pad(`DP4_8),
  .default_value(`default_value)));
ap_DP4_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE)
));
ap_DP4_8_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_8_PINCTRL_0_IE),
  .outen(`DP4_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_8),
  .pad(`DP4_8),
  .default_value(`default_value)));
ap_DP4_8_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP4_8)
));
ap_DP4_8_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_8_OUTFUNC_SEL),
  .gpioouten(`DP4_8_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP4_8_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP4_8),
  .pad_gz(`DP4_8_pad_y)
));
ap_DP4_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_8_PULLEN),
  .pullsel(`DP4_8_PULLSEL),
  .pad_pullup(`DP4_8)
));
ap_DP4_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .pullsel(`DP4_8_PULLSEL)
));
ap_DP4_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_8_PULLEN),
  .pullsel(`DP4_8_PULLSEL),
  .pad_pd(`DP4_8)
));
ap_DP4_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_8),
  .pullen(`DP4_8_PULLEN),
  .pullsel(`DP4_8_PULLSEL)
));
ap_DP4_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD2_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`RGMII1TXD2_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD2_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`RGMII1TXD2_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE)
));
ap_DP4_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_9_PINCTRL_0_IE),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_9),
  .pad(`DP4_9),
  .default_value(`default_value)));
ap_DP4_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE)
));
ap_DP4_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_9_PINCTRL_0_IE),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_9),
  .pad(`DP4_9),
  .default_value(`default_value)));
ap_DP4_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE)
));
ap_DP4_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_9_PINCTRL_0_IE),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_9),
  .pad(`DP4_9),
  .default_value(`default_value)));
ap_DP4_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE)
));
ap_DP4_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_9_PINCTRL_0_IE),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_9),
  .pad(`DP4_9),
  .default_value(`default_value)));
ap_DP4_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE)
));
ap_DP4_9_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_9_PINCTRL_0_IE),
  .outen(`DP4_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_9),
  .pad(`DP4_9),
  .default_value(`default_value)));
ap_DP4_9_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP4_9)
));
ap_DP4_9_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_9_OUTFUNC_SEL),
  .gpioouten(`DP4_9_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP4_9_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP4_9),
  .pad_gz(`DP4_9_pad_y)
));
ap_DP4_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_9_PULLEN),
  .pullsel(`DP4_9_PULLSEL),
  .pad_pullup(`DP4_9)
));
ap_DP4_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .pullsel(`DP4_9_PULLSEL)
));
ap_DP4_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_9_PULLEN),
  .pullsel(`DP4_9_PULLSEL),
  .pad_pd(`DP4_9)
));
ap_DP4_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_9),
  .pullen(`DP4_9_PULLEN),
  .pullsel(`DP4_9_PULLSEL)
));
ap_DP4_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD3_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`RGMII1TXD3_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXD3_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`RGMII1TXD3_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE)
));
ap_DP4_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_10_PINCTRL_0_IE),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_10),
  .pad(`DP4_10),
  .default_value(`default_value)));
ap_DP4_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE)
));
ap_DP4_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_10_PINCTRL_0_IE),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_10),
  .pad(`DP4_10),
  .default_value(`default_value)));
ap_DP4_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE)
));
ap_DP4_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_10_PINCTRL_0_IE),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_10),
  .pad(`DP4_10),
  .default_value(`default_value)));
ap_DP4_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE)
));
ap_DP4_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_10_PINCTRL_0_IE),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_10),
  .pad(`DP4_10),
  .default_value(`default_value)));
ap_DP4_10_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE)
));
ap_DP4_10_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_10_PINCTRL_0_IE),
  .outen(`DP4_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_10),
  .pad(`DP4_10),
  .default_value(`default_value)));
ap_DP4_10_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP4_10)
));
ap_DP4_10_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_10_OUTFUNC_SEL),
  .gpioouten(`DP4_10_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP4_10_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP4_10),
  .pad_gz(`DP4_10_pad_y)
));
ap_DP4_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_10_PULLEN),
  .pullsel(`DP4_10_PULLSEL),
  .pad_pullup(`DP4_10)
));
ap_DP4_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .pullsel(`DP4_10_PULLSEL)
));
ap_DP4_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_10_PULLEN),
  .pullsel(`DP4_10_PULLSEL),
  .pad_pd(`DP4_10)
));
ap_DP4_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_10),
  .pullen(`DP4_10_PULLEN),
  .pullsel(`DP4_10_PULLSEL)
));
ap_DP4_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXCTL_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`RGMII1TXCTL_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1TXCTL_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`RGMII1TXCTL_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE)
));
ap_DP4_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_11_PINCTRL_0_IE),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_11),
  .pad(`DP4_11),
  .default_value(`default_value)));
ap_DP4_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE)
));
ap_DP4_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_11_PINCTRL_0_IE),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_11),
  .pad(`DP4_11),
  .default_value(`default_value)));
ap_DP4_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE)
));
ap_DP4_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_11_PINCTRL_0_IE),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_11),
  .pad(`DP4_11),
  .default_value(`default_value)));
ap_DP4_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE)
));
ap_DP4_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_11_PINCTRL_0_IE),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_11),
  .pad(`DP4_11),
  .default_value(`default_value)));
ap_DP4_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE)
));
ap_DP4_11_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_11_PINCTRL_0_IE),
  .outen(`DP4_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_11),
  .pad(`DP4_11),
  .default_value(`default_value)));
ap_DP4_11_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP4_11)
));
ap_DP4_11_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_11_OUTFUNC_SEL),
  .gpioouten(`DP4_11_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP4_11_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP4_11),
  .pad_gz(`DP4_11_pad_y)
));
ap_DP4_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_11_PULLEN),
  .pullsel(`DP4_11_PULLSEL),
  .pad_pullup(`DP4_11)
));
ap_DP4_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .pullsel(`DP4_11_PULLSEL)
));
ap_DP4_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_11_PULLEN),
  .pullsel(`DP4_11_PULLSEL),
  .pad_pd(`DP4_11)
));
ap_DP4_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_11),
  .pullen(`DP4_11_PULLEN),
  .pullsel(`DP4_11_PULLSEL)
));
ap_DP4_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXCLK_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`RGMII1RXCLK_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXCLK_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`RGMII1RXCLK_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE)
));
ap_DP4_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_12_PINCTRL_0_IE),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_12),
  .pad(`DP4_12),
  .default_value(`default_value)));
ap_DP4_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXCLK_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`FSI4TXCLK_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXCLK_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`FSI4TXCLK_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE)
));
ap_DP4_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_12_PINCTRL_0_IE),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_12),
  .pad(`DP4_12),
  .default_value(`default_value)));
ap_DP4_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE)
));
ap_DP4_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_12_PINCTRL_0_IE),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_12),
  .pad(`DP4_12),
  .default_value(`default_value)));
ap_DP4_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE)
));
ap_DP4_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_12_PINCTRL_0_IE),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_12),
  .pad(`DP4_12),
  .default_value(`default_value)));
ap_DP4_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20B_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`EPWM20B_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE)
));
ap_DP4_12_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_12_PINCTRL_0_IE),
  .outen(`DP4_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_12),
  .pad(`DP4_12),
  .default_value(`default_value)));
ap_DP4_12_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP4_12)
));
ap_DP4_12_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_12_OUTFUNC_SEL),
  .gpioouten(`DP4_12_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP4_12_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP4_12),
  .pad_gz(`DP4_12_pad_y)
));
ap_DP4_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_12_PULLEN),
  .pullsel(`DP4_12_PULLSEL),
  .pad_pullup(`DP4_12)
));
ap_DP4_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .pullsel(`DP4_12_PULLSEL)
));
ap_DP4_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_12_PULLEN),
  .pullsel(`DP4_12_PULLSEL),
  .pad_pd(`DP4_12)
));
ap_DP4_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_12),
  .pullen(`DP4_12_PULLEN),
  .pullsel(`DP4_12_PULLSEL)
));
ap_DP4_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD0_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`RGMII1RXD0_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD0_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`RGMII1RXD0_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE)
));
ap_DP4_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_13_PINCTRL_0_IE),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_13),
  .pad(`DP4_13),
  .default_value(`default_value)));
ap_DP4_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD0_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`FSI4TXD0_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD0_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`FSI4TXD0_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE)
));
ap_DP4_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_13_PINCTRL_0_IE),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_13),
  .pad(`DP4_13),
  .default_value(`default_value)));
ap_DP4_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE)
));
ap_DP4_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_13_PINCTRL_0_IE),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_13),
  .pad(`DP4_13),
  .default_value(`default_value)));
ap_DP4_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE)
));
ap_DP4_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_13_PINCTRL_0_IE),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_13),
  .pad(`DP4_13),
  .default_value(`default_value)));
ap_DP4_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM20A_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`EPWM20A_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE)
));
ap_DP4_13_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_13_PINCTRL_0_IE),
  .outen(`DP4_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_13),
  .pad(`DP4_13),
  .default_value(`default_value)));
ap_DP4_13_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP4_13)
));
ap_DP4_13_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_13_OUTFUNC_SEL),
  .gpioouten(`DP4_13_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP4_13_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP4_13),
  .pad_gz(`DP4_13_pad_y)
));
ap_DP4_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_13_PULLEN),
  .pullsel(`DP4_13_PULLSEL),
  .pad_pullup(`DP4_13)
));
ap_DP4_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .pullsel(`DP4_13_PULLSEL)
));
ap_DP4_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_13_PULLEN),
  .pullsel(`DP4_13_PULLSEL),
  .pad_pd(`DP4_13)
));
ap_DP4_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_13),
  .pullen(`DP4_13_PULLEN),
  .pullsel(`DP4_13_PULLSEL)
));
ap_DP4_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD1_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`RGMII1RXD1_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD1_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`RGMII1RXD1_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE)
));
ap_DP4_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_14_PINCTRL_0_IE),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_14),
  .pad(`DP4_14),
  .default_value(`default_value)));
ap_DP4_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD1_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`FSI4TXD1_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4TXD1_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`FSI4TXD1_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE)
));
ap_DP4_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_14_PINCTRL_0_IE),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_14),
  .pad(`DP4_14),
  .default_value(`default_value)));
ap_DP4_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE)
));
ap_DP4_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_14_PINCTRL_0_IE),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_14),
  .pad(`DP4_14),
  .default_value(`default_value)));
ap_DP4_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE)
));
ap_DP4_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_14_PINCTRL_0_IE),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_14),
  .pad(`DP4_14),
  .default_value(`default_value)));
ap_DP4_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19B_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`EPWM19B_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_14_OUTFUNC_SEL),
  .gpioouten(`DP4_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP4_14_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP4_14),
  .pad_gz(`DP4_14_pad_y)
));
ap_DP4_14_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_14)
));
ap_DP4_14_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE)
));
ap_DP4_14_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_14_PINCTRL_0_IE),
  .outen(`DP4_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_14),
  .pad(`DP4_14),
  .default_value(`default_value)));
ap_DP4_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_14_PULLEN),
  .pullsel(`DP4_14_PULLSEL),
  .pad_pullup(`DP4_14)
));
ap_DP4_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .pullsel(`DP4_14_PULLSEL)
));
ap_DP4_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_14_PULLEN),
  .pullsel(`DP4_14_PULLSEL),
  .pad_pd(`DP4_14)
));
ap_DP4_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_14),
  .pullen(`DP4_14_PULLEN),
  .pullsel(`DP4_14_PULLSEL)
));
ap_DP4_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD2_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`RGMII1RXD2_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD2_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`RGMII1RXD2_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXCLK_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`FSI4RXCLK_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXCLK_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`FSI4RXCLK_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM19A_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`EPWM19A_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_15_OUTFUNC_SEL),
  .gpioouten(`DP4_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`DP4_15_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`DP4_15),
  .pad_gz(`DP4_15_pad_y)
));
ap_DP4_15_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_15)
));
ap_DP4_15_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE)
));
ap_DP4_15_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_15_PINCTRL_0_IE),
  .outen(`DP4_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_15),
  .pad(`DP4_15),
  .default_value(`default_value)));
ap_DP4_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_15_PULLEN),
  .pullsel(`DP4_15_PULLSEL),
  .pad_pullup(`DP4_15)
));
ap_DP4_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .pullsel(`DP4_15_PULLSEL)
));
ap_DP4_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_15_PULLEN),
  .pullsel(`DP4_15_PULLSEL),
  .pad_pd(`DP4_15)
));
ap_DP4_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_15),
  .pullen(`DP4_15_PULLEN),
  .pullsel(`DP4_15_PULLSEL)
));
ap_DP4_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD3_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`RGMII1RXD3_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXD3_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`RGMII1RXD3_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD0_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`FSI4RXD0_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD0_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`FSI4RXD0_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18B_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`EPWM18B_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_16_OUTFUNC_SEL),
  .gpioouten(`DP4_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`DP4_16_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`DP4_16),
  .pad_gz(`DP4_16_pad_y)
));
ap_DP4_16_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_16)
));
ap_DP4_16_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE)
));
ap_DP4_16_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_16_PINCTRL_0_IE),
  .outen(`DP4_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_16),
  .pad(`DP4_16),
  .default_value(`default_value)));
ap_DP4_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_16_PULLEN),
  .pullsel(`DP4_16_PULLSEL),
  .pad_pullup(`DP4_16)
));
ap_DP4_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .pullsel(`DP4_16_PULLSEL)
));
ap_DP4_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_16_PULLEN),
  .pullsel(`DP4_16_PULLSEL),
  .pad_pd(`DP4_16)
));
ap_DP4_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_16),
  .pullen(`DP4_16_PULLEN),
  .pullsel(`DP4_16_PULLSEL)
));
ap_DP4_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXCTL_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`RGMII1RXCTL_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII1RXCTL_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`RGMII1RXCTL_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD1_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`FSI4RXD1_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`FSI4RXD1_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`FSI4RXD1_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM18A_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`EPWM18A_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_17_OUTFUNC_SEL),
  .gpioouten(`DP4_17_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`DP4_17_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`DP4_17),
  .pad_gz(`DP4_17_pad_y)
));
ap_DP4_17_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_17)
));
ap_DP4_17_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE)
));
ap_DP4_17_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_17_PINCTRL_0_IE),
  .outen(`DP4_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_17),
  .pad(`DP4_17),
  .default_value(`default_value)));
ap_DP4_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_17_PULLEN),
  .pullsel(`DP4_17_PULLSEL),
  .pad_pullup(`DP4_17)
));
ap_DP4_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .pullsel(`DP4_17_PULLSEL)
));
ap_DP4_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_17_PULLEN),
  .pullsel(`DP4_17_PULLSEL),
  .pad_pd(`DP4_17)
));
ap_DP4_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_17),
  .pullen(`DP4_17_PULLEN),
  .pullsel(`DP4_17_PULLSEL)
));
ap_DP4_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_18_OUTFUNC_SEL),
  .gpioouten(`DP4_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_18_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_18)
));
ap_DP4_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_18_OUTFUNC_SEL),
  .gpioouten(`DP4_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_18_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_18),
  .pad_gz(`DP4_18_pad_y)
));
ap_DP4_18_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_18_PULLEN),
  .outen(`DP4_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_18)
));
ap_DP4_18_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_18),
  .pullen(`DP4_18_PULLEN),
  .outen(`DP4_18_GPIO_OUTPUT_ENABLE)
));
ap_DP4_18_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_18_PINCTRL_0_IE),
  .outen(`DP4_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_18),
  .pad(`DP4_18),
  .default_value(`default_value)));
ap_DP4_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_18_OUTFUNC_SEL),
  .gpioouten(`DP4_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP4_18_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP4_18)
));
ap_DP4_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_18_OUTFUNC_SEL),
  .gpioouten(`DP4_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17B_OE),
  .od(`DP4_18_PINCTRL_0_OD),
  .func_out(`EPWM17B_OUT),
  .pad(`DP4_18),
  .pad_gz(`DP4_18_pad_y)
));
ap_DP4_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_18_PULLEN),
  .pullsel(`DP4_18_PULLSEL),
  .pad_pullup(`DP4_18)
));
ap_DP4_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_18),
  .pullen(`DP4_18_PULLEN),
  .pullsel(`DP4_18_PULLSEL)
));
ap_DP4_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_18_PULLEN),
  .pullsel(`DP4_18_PULLSEL),
  .pad_pd(`DP4_18)
));
ap_DP4_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_18),
  .pullen(`DP4_18_PULLEN),
  .pullsel(`DP4_18_PULLSEL)
));
ap_DP4_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_19_OUTFUNC_SEL),
  .gpioouten(`DP4_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_19_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_19)
));
ap_DP4_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_19_OUTFUNC_SEL),
  .gpioouten(`DP4_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_19_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_19),
  .pad_gz(`DP4_19_pad_y)
));
ap_DP4_19_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_19_PULLEN),
  .outen(`DP4_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_19)
));
ap_DP4_19_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_19),
  .pullen(`DP4_19_PULLEN),
  .outen(`DP4_19_GPIO_OUTPUT_ENABLE)
));
ap_DP4_19_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_19_PINCTRL_0_IE),
  .outen(`DP4_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_19),
  .pad(`DP4_19),
  .default_value(`default_value)));
ap_DP4_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_19_OUTFUNC_SEL),
  .gpioouten(`DP4_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP4_19_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP4_19)
));
ap_DP4_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_19_OUTFUNC_SEL),
  .gpioouten(`DP4_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM17A_OE),
  .od(`DP4_19_PINCTRL_0_OD),
  .func_out(`EPWM17A_OUT),
  .pad(`DP4_19),
  .pad_gz(`DP4_19_pad_y)
));
ap_DP4_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_19_PULLEN),
  .pullsel(`DP4_19_PULLSEL),
  .pad_pullup(`DP4_19)
));
ap_DP4_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_19),
  .pullen(`DP4_19_PULLEN),
  .pullsel(`DP4_19_PULLSEL)
));
ap_DP4_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_19_PULLEN),
  .pullsel(`DP4_19_PULLSEL),
  .pad_pd(`DP4_19)
));
ap_DP4_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_19),
  .pullen(`DP4_19_PULLEN),
  .pullsel(`DP4_19_PULLSEL)
));
ap_DP4_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`XSPI0CLK_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`XSPI0CLK_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE)
));
ap_DP4_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_20_PINCTRL_0_IE),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_20),
  .pad(`DP4_20),
  .default_value(`default_value)));
ap_DP4_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE)
));
ap_DP4_20_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_20_PINCTRL_0_IE),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_20),
  .pad(`DP4_20),
  .default_value(`default_value)));
ap_DP4_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30A_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`EPWM30A_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0EXTREFCLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MCASP0EXTREFCLK_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE)
));
ap_DP4_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_20_PINCTRL_0_IE),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_20),
  .pad(`DP4_20),
  .default_value(`default_value)));
ap_DP4_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16B_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`EPWM16B_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE)
));
ap_DP4_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_20_PINCTRL_0_IE),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_20),
  .pad(`DP4_20),
  .default_value(`default_value)));
ap_DP4_20_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_20_OUTFUNC_SEL),
  .gpioouten(`DP4_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`DP4_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`DP4_20),
  .pad_gz(`DP4_20_pad_y)
));
ap_DP4_20_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_20)
));
ap_DP4_20_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE)
));
ap_DP4_20_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_20_PINCTRL_0_IE),
  .outen(`DP4_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_20),
  .pad(`DP4_20),
  .default_value(`default_value)));
ap_DP4_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_20_PULLEN),
  .pullsel(`DP4_20_PULLSEL),
  .pad_pullup(`DP4_20)
));
ap_DP4_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .pullsel(`DP4_20_PULLSEL)
));
ap_DP4_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_20_PULLEN),
  .pullsel(`DP4_20_PULLSEL),
  .pad_pd(`DP4_20)
));
ap_DP4_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_20),
  .pullen(`DP4_20_PULLEN),
  .pullsel(`DP4_20_PULLSEL)
));
ap_DP4_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CS0_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`XSPI0CS0_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CS0_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`XSPI0CS0_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE)
));
ap_DP4_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_21_PINCTRL_0_IE),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_21),
  .pad(`DP4_21),
  .default_value(`default_value)));
ap_DP4_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE)
));
ap_DP4_21_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_21_PINCTRL_0_IE),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_21),
  .pad(`DP4_21),
  .default_value(`default_value)));
ap_DP4_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM30B_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`EPWM30B_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKX_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKX_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE)
));
ap_DP4_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_21_PINCTRL_0_IE),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_21),
  .pad(`DP4_21),
  .default_value(`default_value)));
ap_DP4_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM16A_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`EPWM16A_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE)
));
ap_DP4_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_21_PINCTRL_0_IE),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_21),
  .pad(`DP4_21),
  .default_value(`default_value)));
ap_DP4_21_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_21_OUTFUNC_SEL),
  .gpioouten(`DP4_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`DP4_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`DP4_21),
  .pad_gz(`DP4_21_pad_y)
));
ap_DP4_21_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_21)
));
ap_DP4_21_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE)
));
ap_DP4_21_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_21_PINCTRL_0_IE),
  .outen(`DP4_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_21),
  .pad(`DP4_21),
  .default_value(`default_value)));
ap_DP4_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_21_PULLEN),
  .pullsel(`DP4_21_PULLSEL),
  .pad_pullup(`DP4_21)
));
ap_DP4_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .pullsel(`DP4_21_PULLSEL)
));
ap_DP4_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_21_PULLEN),
  .pullsel(`DP4_21_PULLSEL),
  .pad_pd(`DP4_21)
));
ap_DP4_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_21),
  .pullen(`DP4_21_PULLEN),
  .pullsel(`DP4_21_PULLSEL)
));
ap_DP4_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CS1_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`XSPI0CS1_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0CS1_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`XSPI0CS1_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE)
));
ap_DP4_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_22_PINCTRL_0_IE),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_22),
  .pad(`DP4_22),
  .default_value(`default_value)));
ap_DP4_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE)
));
ap_DP4_22_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_22_PINCTRL_0_IE),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_22),
  .pad(`DP4_22),
  .default_value(`default_value)));
ap_DP4_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31A_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`EPWM31A_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSX_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MCASP0AFSX_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE)
));
ap_DP4_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_22_PINCTRL_0_IE),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_22),
  .pad(`DP4_22),
  .default_value(`default_value)));
ap_DP4_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15B_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`EPWM15B_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE)
));
ap_DP4_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_22_PINCTRL_0_IE),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_22),
  .pad(`DP4_22),
  .default_value(`default_value)));
ap_DP4_22_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_22_OUTFUNC_SEL),
  .gpioouten(`DP4_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`DP4_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`DP4_22),
  .pad_gz(`DP4_22_pad_y)
));
ap_DP4_22_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_22)
));
ap_DP4_22_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE)
));
ap_DP4_22_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_22_PINCTRL_0_IE),
  .outen(`DP4_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_22),
  .pad(`DP4_22),
  .default_value(`default_value)));
ap_DP4_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_22_PULLEN),
  .pullsel(`DP4_22_PULLSEL),
  .pad_pullup(`DP4_22)
));
ap_DP4_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .pullsel(`DP4_22_PULLSEL)
));
ap_DP4_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_22_PULLEN),
  .pullsel(`DP4_22_PULLSEL),
  .pad_pd(`DP4_22)
));
ap_DP4_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_22),
  .pullen(`DP4_22_PULLEN),
  .pullsel(`DP4_22_PULLSEL)
));
ap_DP4_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS0_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`XSPI0DS0_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS0_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`XSPI0DS0_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE)
));
ap_DP4_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_23_PINCTRL_0_IE),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_23),
  .pad(`DP4_23),
  .default_value(`default_value)));
ap_DP4_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE)
));
ap_DP4_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_23_PINCTRL_0_IE),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_23),
  .pad(`DP4_23),
  .default_value(`default_value)));
ap_DP4_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM31B_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`EPWM31B_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0ACLKR_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MCASP0ACLKR_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE)
));
ap_DP4_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_23_PINCTRL_0_IE),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_23),
  .pad(`DP4_23),
  .default_value(`default_value)));
ap_DP4_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM15A_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`EPWM15A_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE)
));
ap_DP4_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_23_PINCTRL_0_IE),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_23),
  .pad(`DP4_23),
  .default_value(`default_value)));
ap_DP4_23_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_23_OUTFUNC_SEL),
  .gpioouten(`DP4_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`DP4_23_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`DP4_23),
  .pad_gz(`DP4_23_pad_y)
));
ap_DP4_23_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_23)
));
ap_DP4_23_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE)
));
ap_DP4_23_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_23_PINCTRL_0_IE),
  .outen(`DP4_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_23),
  .pad(`DP4_23),
  .default_value(`default_value)));
ap_DP4_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_23_PULLEN),
  .pullsel(`DP4_23_PULLSEL),
  .pad_pullup(`DP4_23)
));
ap_DP4_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .pullsel(`DP4_23_PULLSEL)
));
ap_DP4_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_23_PULLEN),
  .pullsel(`DP4_23_PULLSEL),
  .pad_pd(`DP4_23)
));
ap_DP4_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_23),
  .pullen(`DP4_23_PULLEN),
  .pullsel(`DP4_23_PULLSEL)
));
ap_DP4_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS1_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`XSPI0DS1_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS1_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`XSPI0DS1_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE)
));
ap_DP4_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_24_PINCTRL_0_IE),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_24),
  .pad(`DP4_24),
  .default_value(`default_value)));
ap_DP4_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE)
));
ap_DP4_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_24_PINCTRL_0_IE),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_24),
  .pad(`DP4_24),
  .default_value(`default_value)));
ap_DP4_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWMSYNCO_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`EPWMSYNCO_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWMSYNCO_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`EPWMSYNCO_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AFSR_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MCASP0AFSR_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE)
));
ap_DP4_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_24_PINCTRL_0_IE),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_24),
  .pad(`DP4_24),
  .default_value(`default_value)));
ap_DP4_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14B_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`EPWM14B_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE)
));
ap_DP4_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_24_PINCTRL_0_IE),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_24),
  .pad(`DP4_24),
  .default_value(`default_value)));
ap_DP4_24_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_24_OUTFUNC_SEL),
  .gpioouten(`DP4_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`DP4_24_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`DP4_24),
  .pad_gz(`DP4_24_pad_y)
));
ap_DP4_24_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_24)
));
ap_DP4_24_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE)
));
ap_DP4_24_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_24_PINCTRL_0_IE),
  .outen(`DP4_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_24),
  .pad(`DP4_24),
  .default_value(`default_value)));
ap_DP4_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_24_PULLEN),
  .pullsel(`DP4_24_PULLSEL),
  .pad_pullup(`DP4_24)
));
ap_DP4_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .pullsel(`DP4_24_PULLSEL)
));
ap_DP4_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_24_PULLEN),
  .pullsel(`DP4_24_PULLSEL),
  .pad_pd(`DP4_24)
));
ap_DP4_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_24),
  .pullen(`DP4_24_PULLEN),
  .pullsel(`DP4_24_PULLSEL)
));
ap_DP4_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS2_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`XSPI0DS2_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS2_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`XSPI0DS2_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE)
));
ap_DP4_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_25_PINCTRL_0_IE),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_25),
  .pad(`DP4_25),
  .default_value(`default_value)));
ap_DP4_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE)
));
ap_DP4_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_25_PINCTRL_0_IE),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_25),
  .pad(`DP4_25),
  .default_value(`default_value)));
ap_DP4_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE)
));
ap_DP4_25_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_25_PINCTRL_0_IE),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_25),
  .pad(`DP4_25),
  .default_value(`default_value)));
ap_DP4_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR0_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`MCASP0AXR0_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE)
));
ap_DP4_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_25_PINCTRL_0_IE),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_25),
  .pad(`DP4_25),
  .default_value(`default_value)));
ap_DP4_25_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM14A_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`EPWM14A_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_25_OUTFUNC_SEL),
  .gpioouten(`DP4_25_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP4_25_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP4_25),
  .pad_gz(`DP4_25_pad_y)
));
ap_DP4_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_25)
));
ap_DP4_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE)
));
ap_DP4_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_25_PINCTRL_0_IE),
  .outen(`DP4_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_25),
  .pad(`DP4_25),
  .default_value(`default_value)));
ap_DP4_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_25_PULLEN),
  .pullsel(`DP4_25_PULLSEL),
  .pad_pullup(`DP4_25)
));
ap_DP4_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .pullsel(`DP4_25_PULLSEL)
));
ap_DP4_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_25_PULLEN),
  .pullsel(`DP4_25_PULLSEL),
  .pad_pd(`DP4_25)
));
ap_DP4_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_25),
  .pullen(`DP4_25_PULLEN),
  .pullsel(`DP4_25_PULLSEL)
));
ap_DP4_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS3_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`XSPI0DS3_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS3_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`XSPI0DS3_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE)
));
ap_DP4_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_26_PINCTRL_0_IE),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_26),
  .pad(`DP4_26),
  .default_value(`default_value)));
ap_DP4_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE)
));
ap_DP4_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_26_PINCTRL_0_IE),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_26),
  .pad(`DP4_26),
  .default_value(`default_value)));
ap_DP4_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE)
));
ap_DP4_26_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_26_PINCTRL_0_IE),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_26),
  .pad(`DP4_26),
  .default_value(`default_value)));
ap_DP4_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR1_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MCASP0AXR1_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE)
));
ap_DP4_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_26_PINCTRL_0_IE),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_26),
  .pad(`DP4_26),
  .default_value(`default_value)));
ap_DP4_26_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13B_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`EPWM13B_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_26_OUTFUNC_SEL),
  .gpioouten(`DP4_26_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP4_26_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP4_26),
  .pad_gz(`DP4_26_pad_y)
));
ap_DP4_26_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_26)
));
ap_DP4_26_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE)
));
ap_DP4_26_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_26_PINCTRL_0_IE),
  .outen(`DP4_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_26),
  .pad(`DP4_26),
  .default_value(`default_value)));
ap_DP4_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_26_PULLEN),
  .pullsel(`DP4_26_PULLSEL),
  .pad_pullup(`DP4_26)
));
ap_DP4_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .pullsel(`DP4_26_PULLSEL)
));
ap_DP4_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_26_PULLEN),
  .pullsel(`DP4_26_PULLSEL),
  .pad_pd(`DP4_26)
));
ap_DP4_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_26),
  .pullen(`DP4_26_PULLEN),
  .pullsel(`DP4_26_PULLSEL)
));
ap_DP4_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS4_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`XSPI0DS4_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS4_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`XSPI0DS4_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE)
));
ap_DP4_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_27_PINCTRL_0_IE),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_27),
  .pad(`DP4_27),
  .default_value(`default_value)));
ap_DP4_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE)
));
ap_DP4_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_27_PINCTRL_0_IE),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_27),
  .pad(`DP4_27),
  .default_value(`default_value)));
ap_DP4_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE)
));
ap_DP4_27_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_27_PINCTRL_0_IE),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_27),
  .pad(`DP4_27),
  .default_value(`default_value)));
ap_DP4_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR2_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`MCASP0AXR2_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE)
));
ap_DP4_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_27_PINCTRL_0_IE),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_27),
  .pad(`DP4_27),
  .default_value(`default_value)));
ap_DP4_27_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM13A_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`EPWM13A_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_27_OUTFUNC_SEL),
  .gpioouten(`DP4_27_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP4_27_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP4_27),
  .pad_gz(`DP4_27_pad_y)
));
ap_DP4_27_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_27)
));
ap_DP4_27_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE)
));
ap_DP4_27_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_27_PINCTRL_0_IE),
  .outen(`DP4_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_27),
  .pad(`DP4_27),
  .default_value(`default_value)));
ap_DP4_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_27_PULLEN),
  .pullsel(`DP4_27_PULLSEL),
  .pad_pullup(`DP4_27)
));
ap_DP4_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .pullsel(`DP4_27_PULLSEL)
));
ap_DP4_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_27_PULLEN),
  .pullsel(`DP4_27_PULLSEL),
  .pad_pd(`DP4_27)
));
ap_DP4_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_27),
  .pullen(`DP4_27_PULLEN),
  .pullsel(`DP4_27_PULLSEL)
));
ap_DP4_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS5_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`XSPI0DS5_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS5_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`XSPI0DS5_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE)
));
ap_DP4_28_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_28_PINCTRL_0_IE),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_28),
  .pad(`DP4_28),
  .default_value(`default_value)));
ap_DP4_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE)
));
ap_DP4_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_28_PINCTRL_0_IE),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_28),
  .pad(`DP4_28),
  .default_value(`default_value)));
ap_DP4_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE)
));
ap_DP4_28_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_28_PINCTRL_0_IE),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_28),
  .pad(`DP4_28),
  .default_value(`default_value)));
ap_DP4_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCASP0AXR3_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`MCASP0AXR3_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE)
));
ap_DP4_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_28_PINCTRL_0_IE),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_28),
  .pad(`DP4_28),
  .default_value(`default_value)));
ap_DP4_28_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12B_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`EPWM12B_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_28_OUTFUNC_SEL),
  .gpioouten(`DP4_28_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP4_28_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP4_28),
  .pad_gz(`DP4_28_pad_y)
));
ap_DP4_28_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_28)
));
ap_DP4_28_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE)
));
ap_DP4_28_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_28_PINCTRL_0_IE),
  .outen(`DP4_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_28),
  .pad(`DP4_28),
  .default_value(`default_value)));
ap_DP4_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_28_PULLEN),
  .pullsel(`DP4_28_PULLSEL),
  .pad_pullup(`DP4_28)
));
ap_DP4_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .pullsel(`DP4_28_PULLSEL)
));
ap_DP4_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_28_PULLEN),
  .pullsel(`DP4_28_PULLSEL),
  .pad_pd(`DP4_28)
));
ap_DP4_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_28),
  .pullen(`DP4_28_PULLEN),
  .pullsel(`DP4_28_PULLSEL)
));
ap_DP4_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS6_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`XSPI0DS6_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS6_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`XSPI0DS6_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE)
));
ap_DP4_29_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_29_PINCTRL_0_IE),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_29),
  .pad(`DP4_29),
  .default_value(`default_value)));
ap_DP4_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE)
));
ap_DP4_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_29_PINCTRL_0_IE),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_29),
  .pad(`DP4_29),
  .default_value(`default_value)));
ap_DP4_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE)
));
ap_DP4_29_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_29_PINCTRL_0_IE),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_29),
  .pad(`DP4_29),
  .default_value(`default_value)));
ap_DP4_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE)
));
ap_DP4_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_29_PINCTRL_0_IE),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_29),
  .pad(`DP4_29),
  .default_value(`default_value)));
ap_DP4_29_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM12A_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`EPWM12A_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_29_OUTFUNC_SEL),
  .gpioouten(`DP4_29_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP4_29_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP4_29),
  .pad_gz(`DP4_29_pad_y)
));
ap_DP4_29_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_29)
));
ap_DP4_29_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE)
));
ap_DP4_29_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_29_PINCTRL_0_IE),
  .outen(`DP4_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_29),
  .pad(`DP4_29),
  .default_value(`default_value)));
ap_DP4_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_29_PULLEN),
  .pullsel(`DP4_29_PULLSEL),
  .pad_pullup(`DP4_29)
));
ap_DP4_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .pullsel(`DP4_29_PULLSEL)
));
ap_DP4_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_29_PULLEN),
  .pullsel(`DP4_29_PULLSEL),
  .pad_pd(`DP4_29)
));
ap_DP4_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_29),
  .pullen(`DP4_29_PULLEN),
  .pullsel(`DP4_29_PULLSEL)
));
ap_DP4_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS7_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`XSPI0DS7_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DS7_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`XSPI0DS7_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11B_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`EPWM11B_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_30_OUTFUNC_SEL),
  .gpioouten(`DP4_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CLK_OE),
  .od(`DP4_30_PINCTRL_0_OD),
  .func_out(`SPI4CLK_OUT),
  .pad(`DP4_30),
  .pad_gz(`DP4_30_pad_y)
));
ap_DP4_30_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_30)
));
ap_DP4_30_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE)
));
ap_DP4_30_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_30_PINCTRL_0_IE),
  .outen(`DP4_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_30),
  .pad(`DP4_30),
  .default_value(`default_value)));
ap_DP4_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_30_PULLEN),
  .pullsel(`DP4_30_PULLSEL),
  .pad_pullup(`DP4_30)
));
ap_DP4_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .pullsel(`DP4_30_PULLSEL)
));
ap_DP4_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_30_PULLEN),
  .pullsel(`DP4_30_PULLSEL),
  .pad_pd(`DP4_30)
));
ap_DP4_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_30),
  .pullen(`DP4_30_PULLEN),
  .pullsel(`DP4_30_PULLSEL)
));
ap_DP4_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DQS_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`XSPI0DQS_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`XSPI0DQS_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`XSPI0DQS_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM11A_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`EPWM11A_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP4_31_OUTFUNC_SEL),
  .gpioouten(`DP4_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4PICO_OE),
  .od(`DP4_31_PINCTRL_0_OD),
  .func_out(`SPI4PICO_OUT),
  .pad(`DP4_31),
  .pad_gz(`DP4_31_pad_y)
));
ap_DP4_31_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP4_31)
));
ap_DP4_31_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE)
));
ap_DP4_31_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP4_31_PINCTRL_0_IE),
  .outen(`DP4_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP4_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP4_31),
  .pad(`DP4_31),
  .default_value(`default_value)));
ap_DP4_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP4_31_PULLEN),
  .pullsel(`DP4_31_PULLSEL),
  .pad_pullup(`DP4_31)
));
ap_DP4_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .pullsel(`DP4_31_PULLSEL)
));
ap_DP4_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP4_31_PULLEN),
  .pullsel(`DP4_31_PULLSEL),
  .pad_pd(`DP4_31)
));
ap_DP4_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP4_31),
  .pullen(`DP4_31_PULLEN),
  .pullsel(`DP4_31_PULLSEL)
));
ap_DP5_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`GMII_MDC_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`GMII_MDC_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`GMII_MDC_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`GMII_MDC_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10B_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`EPWM10B_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_0_OUTFUNC_SEL),
  .gpioouten(`DP5_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4POCI_OE),
  .od(`DP5_0_PINCTRL_0_OD),
  .func_out(`SPI4POCI_OUT),
  .pad(`DP5_0),
  .pad_gz(`DP5_0_pad_y)
));
ap_DP5_0_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_0)
));
ap_DP5_0_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE)
));
ap_DP5_0_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_0_PINCTRL_0_IE),
  .outen(`DP5_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_0),
  .pad(`DP5_0),
  .default_value(`default_value)));
ap_DP5_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_0_PULLEN),
  .pullsel(`DP5_0_PULLSEL),
  .pad_pullup(`DP5_0)
));
ap_DP5_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .pullsel(`DP5_0_PULLSEL)
));
ap_DP5_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_0_PULLEN),
  .pullsel(`DP5_0_PULLSEL),
  .pad_pd(`DP5_0)
));
ap_DP5_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_0),
  .pullen(`DP5_0_PULLEN),
  .pullsel(`DP5_0_PULLSEL)
));
ap_DP5_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`GMII_MDIO_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`GMII_MDIO_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`GMII_MDIO_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`GMII_MDIO_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM10A_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`EPWM10A_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_1_OUTFUNC_SEL),
  .gpioouten(`DP5_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS0_OE),
  .od(`DP5_1_PINCTRL_0_OD),
  .func_out(`SPI4CS0_OUT),
  .pad(`DP5_1),
  .pad_gz(`DP5_1_pad_y)
));
ap_DP5_1_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_1)
));
ap_DP5_1_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE)
));
ap_DP5_1_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_1_PINCTRL_0_IE),
  .outen(`DP5_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_1),
  .pad(`DP5_1),
  .default_value(`default_value)));
ap_DP5_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_1_PULLEN),
  .pullsel(`DP5_1_PULLSEL),
  .pad_pullup(`DP5_1)
));
ap_DP5_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .pullsel(`DP5_1_PULLSEL)
));
ap_DP5_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_1_PULLEN),
  .pullsel(`DP5_1_PULLSEL),
  .pad_pd(`DP5_1)
));
ap_DP5_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_1),
  .pullen(`DP5_1_PULLEN),
  .pullsel(`DP5_1_PULLSEL)
));
ap_DP5_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXCLK_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`RGMII0TXCLK_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXCLK_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`RGMII0TXCLK_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9B_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`EPWM9B_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_2_OUTFUNC_SEL),
  .gpioouten(`DP5_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS1_OE),
  .od(`DP5_2_PINCTRL_0_OD),
  .func_out(`SPI4CS1_OUT),
  .pad(`DP5_2),
  .pad_gz(`DP5_2_pad_y)
));
ap_DP5_2_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_2)
));
ap_DP5_2_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE)
));
ap_DP5_2_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_2_PINCTRL_0_IE),
  .outen(`DP5_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_2),
  .pad(`DP5_2),
  .default_value(`default_value)));
ap_DP5_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_2_PULLEN),
  .pullsel(`DP5_2_PULLSEL),
  .pad_pullup(`DP5_2)
));
ap_DP5_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .pullsel(`DP5_2_PULLSEL)
));
ap_DP5_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_2_PULLEN),
  .pullsel(`DP5_2_PULLSEL),
  .pad_pd(`DP5_2)
));
ap_DP5_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_2),
  .pullen(`DP5_2_PULLEN),
  .pullsel(`DP5_2_PULLSEL)
));
ap_DP5_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD0_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`RGMII0TXD0_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD0_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`RGMII0TXD0_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM9A_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`EPWM9A_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_3_OUTFUNC_SEL),
  .gpioouten(`DP5_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS2_OE),
  .od(`DP5_3_PINCTRL_0_OD),
  .func_out(`SPI4CS2_OUT),
  .pad(`DP5_3),
  .pad_gz(`DP5_3_pad_y)
));
ap_DP5_3_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_3)
));
ap_DP5_3_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE)
));
ap_DP5_3_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_3_PINCTRL_0_IE),
  .outen(`DP5_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_3),
  .pad(`DP5_3),
  .default_value(`default_value)));
ap_DP5_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_3_PULLEN),
  .pullsel(`DP5_3_PULLSEL),
  .pad_pullup(`DP5_3)
));
ap_DP5_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .pullsel(`DP5_3_PULLSEL)
));
ap_DP5_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_3_PULLEN),
  .pullsel(`DP5_3_PULLSEL),
  .pad_pd(`DP5_3)
));
ap_DP5_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_3),
  .pullen(`DP5_3_PULLEN),
  .pullsel(`DP5_3_PULLSEL)
));
ap_DP5_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD1_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`RGMII0TXD1_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD1_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`RGMII0TXD1_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8B_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`EPWM8B_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_4_OUTFUNC_SEL),
  .gpioouten(`DP5_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS3_OE),
  .od(`DP5_4_PINCTRL_0_OD),
  .func_out(`SPI4CS3_OUT),
  .pad(`DP5_4),
  .pad_gz(`DP5_4_pad_y)
));
ap_DP5_4_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_4)
));
ap_DP5_4_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE)
));
ap_DP5_4_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_4_PINCTRL_0_IE),
  .outen(`DP5_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_4),
  .pad(`DP5_4),
  .default_value(`default_value)));
ap_DP5_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_4_PULLEN),
  .pullsel(`DP5_4_PULLSEL),
  .pad_pullup(`DP5_4)
));
ap_DP5_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .pullsel(`DP5_4_PULLSEL)
));
ap_DP5_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_4_PULLEN),
  .pullsel(`DP5_4_PULLSEL),
  .pad_pd(`DP5_4)
));
ap_DP5_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_4),
  .pullen(`DP5_4_PULLEN),
  .pullsel(`DP5_4_PULLSEL)
));
ap_DP5_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD2_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`RGMII0TXD2_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD2_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`RGMII0TXD2_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE)
));
ap_DP5_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_5_PINCTRL_0_IE),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_5),
  .pad(`DP5_5),
  .default_value(`default_value)));
ap_DP5_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE)
));
ap_DP5_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_5_PINCTRL_0_IE),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_5),
  .pad(`DP5_5),
  .default_value(`default_value)));
ap_DP5_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE)
));
ap_DP5_5_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_5_PINCTRL_0_IE),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_5),
  .pad(`DP5_5),
  .default_value(`default_value)));
ap_DP5_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE)
));
ap_DP5_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_5_PINCTRL_0_IE),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_5),
  .pad(`DP5_5),
  .default_value(`default_value)));
ap_DP5_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM8A_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`EPWM8A_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_5_OUTFUNC_SEL),
  .gpioouten(`DP5_5_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`DP5_5_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`DP5_5),
  .pad_gz(`DP5_5_pad_y)
));
ap_DP5_5_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_5)
));
ap_DP5_5_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE)
));
ap_DP5_5_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_5_PINCTRL_0_IE),
  .outen(`DP5_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_5),
  .pad(`DP5_5),
  .default_value(`default_value)));
ap_DP5_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_5_PULLEN),
  .pullsel(`DP5_5_PULLSEL),
  .pad_pullup(`DP5_5)
));
ap_DP5_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .pullsel(`DP5_5_PULLSEL)
));
ap_DP5_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_5_PULLEN),
  .pullsel(`DP5_5_PULLSEL),
  .pad_pd(`DP5_5)
));
ap_DP5_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_5),
  .pullen(`DP5_5_PULLEN),
  .pullsel(`DP5_5_PULLSEL)
));
ap_DP5_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD3_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`RGMII0TXD3_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXD3_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`RGMII0TXD3_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE)
));
ap_DP5_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_6_PINCTRL_0_IE),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_6),
  .pad(`DP5_6),
  .default_value(`default_value)));
ap_DP5_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE)
));
ap_DP5_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_6_PINCTRL_0_IE),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_6),
  .pad(`DP5_6),
  .default_value(`default_value)));
ap_DP5_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE)
));
ap_DP5_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_6_PINCTRL_0_IE),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_6),
  .pad(`DP5_6),
  .default_value(`default_value)));
ap_DP5_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE)
));
ap_DP5_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_6_PINCTRL_0_IE),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_6),
  .pad(`DP5_6),
  .default_value(`default_value)));
ap_DP5_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7B_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`EPWM7B_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_6_OUTFUNC_SEL),
  .gpioouten(`DP5_6_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`DP5_6_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`DP5_6),
  .pad_gz(`DP5_6_pad_y)
));
ap_DP5_6_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_6)
));
ap_DP5_6_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE)
));
ap_DP5_6_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_6_PINCTRL_0_IE),
  .outen(`DP5_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_6),
  .pad(`DP5_6),
  .default_value(`default_value)));
ap_DP5_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_6_PULLEN),
  .pullsel(`DP5_6_PULLSEL),
  .pad_pullup(`DP5_6)
));
ap_DP5_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .pullsel(`DP5_6_PULLSEL)
));
ap_DP5_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_6_PULLEN),
  .pullsel(`DP5_6_PULLSEL),
  .pad_pd(`DP5_6)
));
ap_DP5_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_6),
  .pullen(`DP5_6_PULLEN),
  .pullsel(`DP5_6_PULLSEL)
));
ap_DP5_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXCTL_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`RGMII0TXCTL_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0TXCTL_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`RGMII0TXCTL_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE)
));
ap_DP5_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_7_PINCTRL_0_IE),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_7),
  .pad(`DP5_7),
  .default_value(`default_value)));
ap_DP5_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE)
));
ap_DP5_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_7_PINCTRL_0_IE),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_7),
  .pad(`DP5_7),
  .default_value(`default_value)));
ap_DP5_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE)
));
ap_DP5_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_7_PINCTRL_0_IE),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_7),
  .pad(`DP5_7),
  .default_value(`default_value)));
ap_DP5_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE)
));
ap_DP5_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_7_PINCTRL_0_IE),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_7),
  .pad(`DP5_7),
  .default_value(`default_value)));
ap_DP5_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM7A_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`EPWM7A_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_7_OUTFUNC_SEL),
  .gpioouten(`DP5_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CLK_OE),
  .od(`DP5_7_PINCTRL_0_OD),
  .func_out(`SPI6CLK_OUT),
  .pad(`DP5_7),
  .pad_gz(`DP5_7_pad_y)
));
ap_DP5_7_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_7)
));
ap_DP5_7_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE)
));
ap_DP5_7_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_7_PINCTRL_0_IE),
  .outen(`DP5_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_7),
  .pad(`DP5_7),
  .default_value(`default_value)));
ap_DP5_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_7_PULLEN),
  .pullsel(`DP5_7_PULLSEL),
  .pad_pullup(`DP5_7)
));
ap_DP5_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .pullsel(`DP5_7_PULLSEL)
));
ap_DP5_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_7_PULLEN),
  .pullsel(`DP5_7_PULLSEL),
  .pad_pd(`DP5_7)
));
ap_DP5_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_7),
  .pullen(`DP5_7_PULLEN),
  .pullsel(`DP5_7_PULLSEL)
));
ap_DP5_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXCLK_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`RGMII0RXCLK_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXCLK_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`RGMII0RXCLK_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE)
));
ap_DP5_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_8_PINCTRL_0_IE),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_8),
  .pad(`DP5_8),
  .default_value(`default_value)));
ap_DP5_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE)
));
ap_DP5_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_8_PINCTRL_0_IE),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_8),
  .pad(`DP5_8),
  .default_value(`default_value)));
ap_DP5_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE)
));
ap_DP5_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_8_PINCTRL_0_IE),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_8),
  .pad(`DP5_8),
  .default_value(`default_value)));
ap_DP5_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE)
));
ap_DP5_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_8_PINCTRL_0_IE),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_8),
  .pad(`DP5_8),
  .default_value(`default_value)));
ap_DP5_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6B_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`EPWM6B_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_8_OUTFUNC_SEL),
  .gpioouten(`DP5_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6PICO_OE),
  .od(`DP5_8_PINCTRL_0_OD),
  .func_out(`SPI6PICO_OUT),
  .pad(`DP5_8),
  .pad_gz(`DP5_8_pad_y)
));
ap_DP5_8_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_8)
));
ap_DP5_8_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE)
));
ap_DP5_8_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_8_PINCTRL_0_IE),
  .outen(`DP5_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_8),
  .pad(`DP5_8),
  .default_value(`default_value)));
ap_DP5_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_8_PULLEN),
  .pullsel(`DP5_8_PULLSEL),
  .pad_pullup(`DP5_8)
));
ap_DP5_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .pullsel(`DP5_8_PULLSEL)
));
ap_DP5_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_8_PULLEN),
  .pullsel(`DP5_8_PULLSEL),
  .pad_pd(`DP5_8)
));
ap_DP5_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_8),
  .pullen(`DP5_8_PULLEN),
  .pullsel(`DP5_8_PULLSEL)
));
ap_DP5_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD0_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`RGMII0RXD0_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD0_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`RGMII0RXD0_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE)
));
ap_DP5_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_9_PINCTRL_0_IE),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_9),
  .pad(`DP5_9),
  .default_value(`default_value)));
ap_DP5_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CLK_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`MIBSPI0CLK_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE)
));
ap_DP5_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_9_PINCTRL_0_IE),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_9),
  .pad(`DP5_9),
  .default_value(`default_value)));
ap_DP5_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE)
));
ap_DP5_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_9_PINCTRL_0_IE),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_9),
  .pad(`DP5_9),
  .default_value(`default_value)));
ap_DP5_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE)
));
ap_DP5_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_9_PINCTRL_0_IE),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_9),
  .pad(`DP5_9),
  .default_value(`default_value)));
ap_DP5_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM6A_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`EPWM6A_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_9_OUTFUNC_SEL),
  .gpioouten(`DP5_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6POCI_OE),
  .od(`DP5_9_PINCTRL_0_OD),
  .func_out(`SPI6POCI_OUT),
  .pad(`DP5_9),
  .pad_gz(`DP5_9_pad_y)
));
ap_DP5_9_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_9)
));
ap_DP5_9_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE)
));
ap_DP5_9_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_9_PINCTRL_0_IE),
  .outen(`DP5_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_9),
  .pad(`DP5_9),
  .default_value(`default_value)));
ap_DP5_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_9_PULLEN),
  .pullsel(`DP5_9_PULLSEL),
  .pad_pullup(`DP5_9)
));
ap_DP5_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .pullsel(`DP5_9_PULLSEL)
));
ap_DP5_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_9_PULLEN),
  .pullsel(`DP5_9_PULLSEL),
  .pad_pd(`DP5_9)
));
ap_DP5_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_9),
  .pullen(`DP5_9_PULLEN),
  .pullsel(`DP5_9_PULLSEL)
));
ap_DP5_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD1_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`RGMII0RXD1_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD1_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`RGMII0RXD1_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE)
));
ap_DP5_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_10_PINCTRL_0_IE),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_10),
  .pad(`DP5_10),
  .default_value(`default_value)));
ap_DP5_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0PICO_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`MIBSPI0PICO_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE)
));
ap_DP5_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_10_PINCTRL_0_IE),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_10),
  .pad(`DP5_10),
  .default_value(`default_value)));
ap_DP5_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE)
));
ap_DP5_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_10_PINCTRL_0_IE),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_10),
  .pad(`DP5_10),
  .default_value(`default_value)));
ap_DP5_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE)
));
ap_DP5_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_10_PINCTRL_0_IE),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_10),
  .pad(`DP5_10),
  .default_value(`default_value)));
ap_DP5_10_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5B_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`EPWM5B_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_10_OUTFUNC_SEL),
  .gpioouten(`DP5_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS0_OE),
  .od(`DP5_10_PINCTRL_0_OD),
  .func_out(`SPI6CS0_OUT),
  .pad(`DP5_10),
  .pad_gz(`DP5_10_pad_y)
));
ap_DP5_10_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_10)
));
ap_DP5_10_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE)
));
ap_DP5_10_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_10_PINCTRL_0_IE),
  .outen(`DP5_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_10),
  .pad(`DP5_10),
  .default_value(`default_value)));
ap_DP5_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_10_PULLEN),
  .pullsel(`DP5_10_PULLSEL),
  .pad_pullup(`DP5_10)
));
ap_DP5_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .pullsel(`DP5_10_PULLSEL)
));
ap_DP5_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_10_PULLEN),
  .pullsel(`DP5_10_PULLSEL),
  .pad_pd(`DP5_10)
));
ap_DP5_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_10),
  .pullen(`DP5_10_PULLEN),
  .pullsel(`DP5_10_PULLSEL)
));
ap_DP5_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD2_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`RGMII0RXD2_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD2_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`RGMII0RXD2_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE)
));
ap_DP5_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_11_PINCTRL_0_IE),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_11),
  .pad(`DP5_11),
  .default_value(`default_value)));
ap_DP5_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0POCI_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`MIBSPI0POCI_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE)
));
ap_DP5_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_11_PINCTRL_0_IE),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_11),
  .pad(`DP5_11),
  .default_value(`default_value)));
ap_DP5_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE)
));
ap_DP5_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_11_PINCTRL_0_IE),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_11),
  .pad(`DP5_11),
  .default_value(`default_value)));
ap_DP5_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE)
));
ap_DP5_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_11_PINCTRL_0_IE),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_11),
  .pad(`DP5_11),
  .default_value(`default_value)));
ap_DP5_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM5A_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`EPWM5A_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_11_OUTFUNC_SEL),
  .gpioouten(`DP5_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS1_OE),
  .od(`DP5_11_PINCTRL_0_OD),
  .func_out(`SPI6CS1_OUT),
  .pad(`DP5_11),
  .pad_gz(`DP5_11_pad_y)
));
ap_DP5_11_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_11)
));
ap_DP5_11_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE)
));
ap_DP5_11_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_11_PINCTRL_0_IE),
  .outen(`DP5_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_11),
  .pad(`DP5_11),
  .default_value(`default_value)));
ap_DP5_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_11_PULLEN),
  .pullsel(`DP5_11_PULLSEL),
  .pad_pullup(`DP5_11)
));
ap_DP5_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .pullsel(`DP5_11_PULLSEL)
));
ap_DP5_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_11_PULLEN),
  .pullsel(`DP5_11_PULLSEL),
  .pad_pd(`DP5_11)
));
ap_DP5_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_11),
  .pullen(`DP5_11_PULLEN),
  .pullsel(`DP5_11_PULLSEL)
));
ap_DP5_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD3_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`RGMII0RXD3_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXD3_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`RGMII0RXD3_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE)
));
ap_DP5_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_12_PINCTRL_0_IE),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_12),
  .pad(`DP5_12),
  .default_value(`default_value)));
ap_DP5_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE)
));
ap_DP5_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_12_PINCTRL_0_IE),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_12),
  .pad(`DP5_12),
  .default_value(`default_value)));
ap_DP5_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE)
));
ap_DP5_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_12_PINCTRL_0_IE),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_12),
  .pad(`DP5_12),
  .default_value(`default_value)));
ap_DP5_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE)
));
ap_DP5_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_12_PINCTRL_0_IE),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_12),
  .pad(`DP5_12),
  .default_value(`default_value)));
ap_DP5_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4B_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`EPWM4B_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_12_OUTFUNC_SEL),
  .gpioouten(`DP5_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS2_OE),
  .od(`DP5_12_PINCTRL_0_OD),
  .func_out(`SPI6CS2_OUT),
  .pad(`DP5_12),
  .pad_gz(`DP5_12_pad_y)
));
ap_DP5_12_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_12)
));
ap_DP5_12_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE)
));
ap_DP5_12_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_12_PINCTRL_0_IE),
  .outen(`DP5_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_12),
  .pad(`DP5_12),
  .default_value(`default_value)));
ap_DP5_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_12_PULLEN),
  .pullsel(`DP5_12_PULLSEL),
  .pad_pullup(`DP5_12)
));
ap_DP5_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .pullsel(`DP5_12_PULLSEL)
));
ap_DP5_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_12_PULLEN),
  .pullsel(`DP5_12_PULLSEL),
  .pad_pd(`DP5_12)
));
ap_DP5_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_12),
  .pullen(`DP5_12_PULLEN),
  .pullsel(`DP5_12_PULLSEL)
));
ap_DP5_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXCTL_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`RGMII0RXCTL_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII0RXCTL_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`RGMII0RXCTL_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE)
));
ap_DP5_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_13_PINCTRL_0_IE),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_13),
  .pad(`DP5_13),
  .default_value(`default_value)));
ap_DP5_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE)
));
ap_DP5_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_13_PINCTRL_0_IE),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_13),
  .pad(`DP5_13),
  .default_value(`default_value)));
ap_DP5_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE)
));
ap_DP5_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_13_PINCTRL_0_IE),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_13),
  .pad(`DP5_13),
  .default_value(`default_value)));
ap_DP5_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE)
));
ap_DP5_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_13_PINCTRL_0_IE),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_13),
  .pad(`DP5_13),
  .default_value(`default_value)));
ap_DP5_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM4A_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`EPWM4A_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_13_OUTFUNC_SEL),
  .gpioouten(`DP5_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS3_OE),
  .od(`DP5_13_PINCTRL_0_OD),
  .func_out(`SPI6CS3_OUT),
  .pad(`DP5_13),
  .pad_gz(`DP5_13_pad_y)
));
ap_DP5_13_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_13)
));
ap_DP5_13_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE)
));
ap_DP5_13_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_13_PINCTRL_0_IE),
  .outen(`DP5_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_13),
  .pad(`DP5_13),
  .default_value(`default_value)));
ap_DP5_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_13_PULLEN),
  .pullsel(`DP5_13_PULLSEL),
  .pad_pullup(`DP5_13)
));
ap_DP5_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .pullsel(`DP5_13_PULLSEL)
));
ap_DP5_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_13_PULLEN),
  .pullsel(`DP5_13_PULLSEL),
  .pad_pd(`DP5_13)
));
ap_DP5_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_13),
  .pullen(`DP5_13_PULLEN),
  .pullsel(`DP5_13_PULLSEL)
));
ap_DP5_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCLK_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`TPIUCLK_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCLK_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`TPIUCLK_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE)
));
ap_DP5_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_14_PINCTRL_0_IE),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_14),
  .pad(`DP5_14),
  .default_value(`default_value)));
ap_DP5_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE)
));
ap_DP5_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_14_PINCTRL_0_IE),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_14),
  .pad(`DP5_14),
  .default_value(`default_value)));
ap_DP5_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0A_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`MCPWM0A_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE)
));
ap_DP5_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_14_PINCTRL_0_IE),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_14),
  .pad(`DP5_14),
  .default_value(`default_value)));
ap_DP5_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_14_OUTFUNC_SEL),
  .gpioouten(`DP5_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CLK_OE),
  .od(`DP5_14_PINCTRL_0_OD),
  .func_out(`SPI7CLK_OUT),
  .pad(`DP5_14),
  .pad_gz(`DP5_14_pad_y)
));
ap_DP5_14_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_14)
));
ap_DP5_14_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE)
));
ap_DP5_14_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_14_PINCTRL_0_IE),
  .outen(`DP5_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_14),
  .pad(`DP5_14),
  .default_value(`default_value)));
ap_DP5_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_14_PULLEN),
  .pullsel(`DP5_14_PULLSEL),
  .pad_pullup(`DP5_14)
));
ap_DP5_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .pullsel(`DP5_14_PULLSEL)
));
ap_DP5_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_14_PULLEN),
  .pullsel(`DP5_14_PULLSEL),
  .pad_pd(`DP5_14)
));
ap_DP5_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_14),
  .pullen(`DP5_14_PULLEN),
  .pullsel(`DP5_14_PULLSEL)
));
ap_DP5_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCTL_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`TPIUCTL_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUCTL_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`TPIUCTL_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE)
));
ap_DP5_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_15_PINCTRL_0_IE),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_15),
  .pad(`DP5_15),
  .default_value(`default_value)));
ap_DP5_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE)
));
ap_DP5_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_15_PINCTRL_0_IE),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_15),
  .pad(`DP5_15),
  .default_value(`default_value)));
ap_DP5_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0B_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`MCPWM0B_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE)
));
ap_DP5_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_15_PINCTRL_0_IE),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_15),
  .pad(`DP5_15),
  .default_value(`default_value)));
ap_DP5_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_15_OUTFUNC_SEL),
  .gpioouten(`DP5_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7PICO_OE),
  .od(`DP5_15_PINCTRL_0_OD),
  .func_out(`SPI7PICO_OUT),
  .pad(`DP5_15),
  .pad_gz(`DP5_15_pad_y)
));
ap_DP5_15_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_15)
));
ap_DP5_15_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE)
));
ap_DP5_15_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_15_PINCTRL_0_IE),
  .outen(`DP5_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_15),
  .pad(`DP5_15),
  .default_value(`default_value)));
ap_DP5_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_15_PULLEN),
  .pullsel(`DP5_15_PULLSEL),
  .pad_pullup(`DP5_15)
));
ap_DP5_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .pullsel(`DP5_15_PULLSEL)
));
ap_DP5_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_15_PULLEN),
  .pullsel(`DP5_15_PULLSEL),
  .pad_pd(`DP5_15)
));
ap_DP5_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_15),
  .pullen(`DP5_15_PULLEN),
  .pullsel(`DP5_15_PULLSEL)
));
ap_DP5_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA0_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`TPIUDATA0_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA0_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`TPIUDATA0_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE)
));
ap_DP5_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_16_PINCTRL_0_IE),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_16),
  .pad(`DP5_16),
  .default_value(`default_value)));
ap_DP5_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE)
));
ap_DP5_16_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_16_PINCTRL_0_IE),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_16),
  .pad(`DP5_16),
  .default_value(`default_value)));
ap_DP5_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0C_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`MCPWM0C_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE)
));
ap_DP5_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_16_PINCTRL_0_IE),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_16),
  .pad(`DP5_16),
  .default_value(`default_value)));
ap_DP5_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_16_OUTFUNC_SEL),
  .gpioouten(`DP5_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7POCI_OE),
  .od(`DP5_16_PINCTRL_0_OD),
  .func_out(`SPI7POCI_OUT),
  .pad(`DP5_16),
  .pad_gz(`DP5_16_pad_y)
));
ap_DP5_16_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_16)
));
ap_DP5_16_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE)
));
ap_DP5_16_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_16_PINCTRL_0_IE),
  .outen(`DP5_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_16),
  .pad(`DP5_16),
  .default_value(`default_value)));
ap_DP5_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_16_PULLEN),
  .pullsel(`DP5_16_PULLSEL),
  .pad_pullup(`DP5_16)
));
ap_DP5_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .pullsel(`DP5_16_PULLSEL)
));
ap_DP5_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_16_PULLEN),
  .pullsel(`DP5_16_PULLSEL),
  .pad_pd(`DP5_16)
));
ap_DP5_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_16),
  .pullen(`DP5_16_PULLEN),
  .pullsel(`DP5_16_PULLSEL)
));
ap_DP5_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA1_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`TPIUDATA1_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA1_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`TPIUDATA1_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE)
));
ap_DP5_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_17_PINCTRL_0_IE),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_17),
  .pad(`DP5_17),
  .default_value(`default_value)));
ap_DP5_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE)
));
ap_DP5_17_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_17_PINCTRL_0_IE),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_17),
  .pad(`DP5_17),
  .default_value(`default_value)));
ap_DP5_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0D_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`MCPWM0D_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE)
));
ap_DP5_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_17_PINCTRL_0_IE),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_17),
  .pad(`DP5_17),
  .default_value(`default_value)));
ap_DP5_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_17_OUTFUNC_SEL),
  .gpioouten(`DP5_17_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS0_OE),
  .od(`DP5_17_PINCTRL_0_OD),
  .func_out(`SPI7CS0_OUT),
  .pad(`DP5_17),
  .pad_gz(`DP5_17_pad_y)
));
ap_DP5_17_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_17)
));
ap_DP5_17_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE)
));
ap_DP5_17_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_17_PINCTRL_0_IE),
  .outen(`DP5_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_17),
  .pad(`DP5_17),
  .default_value(`default_value)));
ap_DP5_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_17_PULLEN),
  .pullsel(`DP5_17_PULLSEL),
  .pad_pullup(`DP5_17)
));
ap_DP5_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .pullsel(`DP5_17_PULLSEL)
));
ap_DP5_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_17_PULLEN),
  .pullsel(`DP5_17_PULLSEL),
  .pad_pd(`DP5_17)
));
ap_DP5_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_17),
  .pullen(`DP5_17_PULLEN),
  .pullsel(`DP5_17_PULLSEL)
));
ap_DP5_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA2_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`TPIUDATA2_OUT),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA2_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`TPIUDATA2_OUT),
  .pad(`DP5_18),
  .pad_gz(`DP5_18_pad_y)
));
ap_DP5_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP5_18),
  .pad_gz(`DP5_18_pad_y)
));
ap_DP5_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_18),
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE)
));
ap_DP5_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_18_PINCTRL_0_IE),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_18),
  .pad(`DP5_18),
  .default_value(`default_value)));
ap_DP5_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0E_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`MCPWM0E_OUT),
  .pad(`DP5_18),
  .pad_gz(`DP5_18_pad_y)
));
ap_DP5_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_18),
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE)
));
ap_DP5_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_18_PINCTRL_0_IE),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_18),
  .pad(`DP5_18),
  .default_value(`default_value)));
ap_DP5_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP5_18),
  .pad_gz(`DP5_18_pad_y)
));
ap_DP5_18_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_18_OUTFUNC_SEL),
  .gpioouten(`DP5_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS1_OE),
  .od(`DP5_18_PINCTRL_0_OD),
  .func_out(`SPI7CS1_OUT),
  .pad(`DP5_18),
  .pad_gz(`DP5_18_pad_y)
));
ap_DP5_18_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_18)
));
ap_DP5_18_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_18),
  .pullen(`DP5_18_PULLEN),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE)
));
ap_DP5_18_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_18_PINCTRL_0_IE),
  .outen(`DP5_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_18),
  .pad(`DP5_18),
  .default_value(`default_value)));
ap_DP5_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_18_PULLEN),
  .pullsel(`DP5_18_PULLSEL),
  .pad_pullup(`DP5_18)
));
ap_DP5_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_18),
  .pullen(`DP5_18_PULLEN),
  .pullsel(`DP5_18_PULLSEL)
));
ap_DP5_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_18_PULLEN),
  .pullsel(`DP5_18_PULLSEL),
  .pad_pd(`DP5_18)
));
ap_DP5_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_18),
  .pullen(`DP5_18_PULLEN),
  .pullsel(`DP5_18_PULLSEL)
));
ap_DP5_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA3_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`TPIUDATA3_OUT),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`TPIUDATA3_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`TPIUDATA3_OUT),
  .pad(`DP5_19),
  .pad_gz(`DP5_19_pad_y)
));
ap_DP5_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP5_19),
  .pad_gz(`DP5_19_pad_y)
));
ap_DP5_19_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_19),
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE)
));
ap_DP5_19_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_19_PINCTRL_0_IE),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_19),
  .pad(`DP5_19),
  .default_value(`default_value)));
ap_DP5_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM0F_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`MCPWM0F_OUT),
  .pad(`DP5_19),
  .pad_gz(`DP5_19_pad_y)
));
ap_DP5_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_19),
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE)
));
ap_DP5_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_19_PINCTRL_0_IE),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_19),
  .pad(`DP5_19),
  .default_value(`default_value)));
ap_DP5_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP5_19),
  .pad_gz(`DP5_19_pad_y)
));
ap_DP5_19_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_19_OUTFUNC_SEL),
  .gpioouten(`DP5_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS2_OE),
  .od(`DP5_19_PINCTRL_0_OD),
  .func_out(`SPI7CS2_OUT),
  .pad(`DP5_19),
  .pad_gz(`DP5_19_pad_y)
));
ap_DP5_19_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_19)
));
ap_DP5_19_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_19),
  .pullen(`DP5_19_PULLEN),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE)
));
ap_DP5_19_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_19_PINCTRL_0_IE),
  .outen(`DP5_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_19),
  .pad(`DP5_19),
  .default_value(`default_value)));
ap_DP5_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_19_PULLEN),
  .pullsel(`DP5_19_PULLSEL),
  .pad_pullup(`DP5_19)
));
ap_DP5_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_19),
  .pullen(`DP5_19_PULLEN),
  .pullsel(`DP5_19_PULLSEL)
));
ap_DP5_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_19_PULLEN),
  .pullsel(`DP5_19_PULLSEL),
  .pad_pd(`DP5_19)
));
ap_DP5_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_19),
  .pullen(`DP5_19_PULLEN),
  .pullsel(`DP5_19_PULLSEL)
));
ap_DP5_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CLK_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`SPI2CLK_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE)
));
ap_DP5_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_20_PINCTRL_0_IE),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_20),
  .pad(`DP5_20),
  .default_value(`default_value)));
ap_DP5_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE)
));
ap_DP5_20_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_20_PINCTRL_0_IE),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_20),
  .pad(`DP5_20),
  .default_value(`default_value)));
ap_DP5_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL0_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL0_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1A_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`MCPWM1A_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE)
));
ap_DP5_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_20_PINCTRL_0_IE),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_20),
  .pad(`DP5_20),
  .default_value(`default_value)));
ap_DP5_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0B_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`EPWM0B_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_20_OUTFUNC_SEL),
  .gpioouten(`DP5_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS3_OE),
  .od(`DP5_20_PINCTRL_0_OD),
  .func_out(`SPI7CS3_OUT),
  .pad(`DP5_20),
  .pad_gz(`DP5_20_pad_y)
));
ap_DP5_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_20)
));
ap_DP5_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE)
));
ap_DP5_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_20_PINCTRL_0_IE),
  .outen(`DP5_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_20),
  .pad(`DP5_20),
  .default_value(`default_value)));
ap_DP5_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_20_PULLEN),
  .pullsel(`DP5_20_PULLSEL),
  .pad_pullup(`DP5_20)
));
ap_DP5_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .pullsel(`DP5_20_PULLSEL)
));
ap_DP5_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_20_PULLEN),
  .pullsel(`DP5_20_PULLSEL),
  .pad_pd(`DP5_20)
));
ap_DP5_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_20),
  .pullen(`DP5_20_PULLEN),
  .pullsel(`DP5_20_PULLSEL)
));
ap_DP5_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2PICO_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`SPI2PICO_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE)
));
ap_DP5_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_21_PINCTRL_0_IE),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_21),
  .pad(`DP5_21),
  .default_value(`default_value)));
ap_DP5_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE)
));
ap_DP5_21_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_21_PINCTRL_0_IE),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_21),
  .pad(`DP5_21),
  .default_value(`default_value)));
ap_DP5_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL1_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL1_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1B_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`MCPWM1B_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE)
));
ap_DP5_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_21_PINCTRL_0_IE),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_21),
  .pad(`DP5_21),
  .default_value(`default_value)));
ap_DP5_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_21_OUTFUNC_SEL),
  .gpioouten(`DP5_21_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP5_21_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP5_21),
  .pad_gz(`DP5_21_pad_y)
));
ap_DP5_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_21)
));
ap_DP5_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE)
));
ap_DP5_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_21_PINCTRL_0_IE),
  .outen(`DP5_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_21),
  .pad(`DP5_21),
  .default_value(`default_value)));
ap_DP5_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_21_PULLEN),
  .pullsel(`DP5_21_PULLSEL),
  .pad_pullup(`DP5_21)
));
ap_DP5_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .pullsel(`DP5_21_PULLSEL)
));
ap_DP5_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_21_PULLEN),
  .pullsel(`DP5_21_PULLSEL),
  .pad_pd(`DP5_21)
));
ap_DP5_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_21),
  .pullen(`DP5_21_PULLEN),
  .pullsel(`DP5_21_PULLSEL)
));
ap_DP5_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2POCI_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`SPI2POCI_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE)
));
ap_DP5_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_22_PINCTRL_0_IE),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_22),
  .pad(`DP5_22),
  .default_value(`default_value)));
ap_DP5_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE)
));
ap_DP5_22_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_22_PINCTRL_0_IE),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_22),
  .pad(`DP5_22),
  .default_value(`default_value)));
ap_DP5_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL0_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL0_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1C_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`MCPWM1C_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE)
));
ap_DP5_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_22_PINCTRL_0_IE),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_22),
  .pad(`DP5_22),
  .default_value(`default_value)));
ap_DP5_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM0A_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`EPWM0A_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_22_OUTFUNC_SEL),
  .gpioouten(`DP5_22_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP5_22_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP5_22),
  .pad_gz(`DP5_22_pad_y)
));
ap_DP5_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_22)
));
ap_DP5_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE)
));
ap_DP5_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_22_PINCTRL_0_IE),
  .outen(`DP5_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_22),
  .pad(`DP5_22),
  .default_value(`default_value)));
ap_DP5_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_22_PULLEN),
  .pullsel(`DP5_22_PULLSEL),
  .pad_pullup(`DP5_22)
));
ap_DP5_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .pullsel(`DP5_22_PULLSEL)
));
ap_DP5_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_22_PULLEN),
  .pullsel(`DP5_22_PULLSEL),
  .pad_pd(`DP5_22)
));
ap_DP5_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_22),
  .pullen(`DP5_22_PULLEN),
  .pullsel(`DP5_22_PULLSEL)
));
ap_DP5_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS0_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`SPI2CS0_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE)
));
ap_DP5_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_23_PINCTRL_0_IE),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_23),
  .pad(`DP5_23),
  .default_value(`default_value)));
ap_DP5_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE)
));
ap_DP5_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_23_PINCTRL_0_IE),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_23),
  .pad(`DP5_23),
  .default_value(`default_value)));
ap_DP5_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL1_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL1_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1D_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`MCPWM1D_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE)
));
ap_DP5_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_23_PINCTRL_0_IE),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_23),
  .pad(`DP5_23),
  .default_value(`default_value)));
ap_DP5_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE)
));
ap_DP5_23_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_23_PINCTRL_0_IE),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_23),
  .pad(`DP5_23),
  .default_value(`default_value)));
ap_DP5_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_23_OUTFUNC_SEL),
  .gpioouten(`DP5_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS1_OE),
  .od(`DP5_23_PINCTRL_0_OD),
  .func_out(`SPI5CS1_OUT),
  .pad(`DP5_23),
  .pad_gz(`DP5_23_pad_y)
));
ap_DP5_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_23)
));
ap_DP5_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE)
));
ap_DP5_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_23_PINCTRL_0_IE),
  .outen(`DP5_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_23),
  .pad(`DP5_23),
  .default_value(`default_value)));
ap_DP5_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_23_PULLEN),
  .pullsel(`DP5_23_PULLSEL),
  .pad_pullup(`DP5_23)
));
ap_DP5_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .pullsel(`DP5_23_PULLSEL)
));
ap_DP5_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_23_PULLEN),
  .pullsel(`DP5_23_PULLSEL),
  .pad_pd(`DP5_23)
));
ap_DP5_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_23),
  .pullen(`DP5_23_PULLEN),
  .pullsel(`DP5_23_PULLSEL)
));
ap_DP5_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE)
));
ap_DP5_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_24_PINCTRL_0_IE),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_24),
  .pad(`DP5_24),
  .default_value(`default_value)));
ap_DP5_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS1_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`SPI2CS1_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE)
));
ap_DP5_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_24_PINCTRL_0_IE),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_24),
  .pad(`DP5_24),
  .default_value(`default_value)));
ap_DP5_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL2_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL2_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1E_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`MCPWM1E_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE)
));
ap_DP5_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_24_PINCTRL_0_IE),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_24),
  .pad(`DP5_24),
  .default_value(`default_value)));
ap_DP5_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE)
));
ap_DP5_24_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_24_PINCTRL_0_IE),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_24),
  .pad(`DP5_24),
  .default_value(`default_value)));
ap_DP5_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_24_OUTFUNC_SEL),
  .gpioouten(`DP5_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS2_OE),
  .od(`DP5_24_PINCTRL_0_OD),
  .func_out(`SPI5CS2_OUT),
  .pad(`DP5_24),
  .pad_gz(`DP5_24_pad_y)
));
ap_DP5_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_24)
));
ap_DP5_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE)
));
ap_DP5_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_24_PINCTRL_0_IE),
  .outen(`DP5_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_24),
  .pad(`DP5_24),
  .default_value(`default_value)));
ap_DP5_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_24_PULLEN),
  .pullsel(`DP5_24_PULLSEL),
  .pad_pullup(`DP5_24)
));
ap_DP5_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .pullsel(`DP5_24_PULLSEL)
));
ap_DP5_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_24_PULLEN),
  .pullsel(`DP5_24_PULLSEL),
  .pad_pd(`DP5_24)
));
ap_DP5_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_24),
  .pullen(`DP5_24_PULLEN),
  .pullsel(`DP5_24_PULLSEL)
));
ap_DP5_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP5_25),
  .pad_gz(`DP5_25_pad_y)
));
ap_DP5_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE)
));
ap_DP5_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_25_PINCTRL_0_IE),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_25),
  .pad(`DP5_25),
  .default_value(`default_value)));
ap_DP5_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS2_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`SPI2CS2_OUT),
  .pad(`DP5_25),
  .pad_gz(`DP5_25_pad_y)
));
ap_DP5_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE)
));
ap_DP5_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_25_PINCTRL_0_IE),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_25),
  .pad(`DP5_25),
  .default_value(`default_value)));
ap_DP5_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`ADC7EXTMUXSEL3_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`ADC7EXTMUXSEL3_OUT),
  .pad(`DP5_25),
  .pad_gz(`DP5_25_pad_y)
));
ap_DP5_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM1F_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`MCPWM1F_OUT),
  .pad(`DP5_25),
  .pad_gz(`DP5_25_pad_y)
));
ap_DP5_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE)
));
ap_DP5_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_25_PINCTRL_0_IE),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_25),
  .pad(`DP5_25),
  .default_value(`default_value)));
ap_DP5_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_25_OUTFUNC_SEL),
  .gpioouten(`DP5_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS3_OE),
  .od(`DP5_25_PINCTRL_0_OD),
  .func_out(`SPI5CS3_OUT),
  .pad(`DP5_25),
  .pad_gz(`DP5_25_pad_y)
));
ap_DP5_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_25)
));
ap_DP5_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE)
));
ap_DP5_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP5_25_PINCTRL_0_IE),
  .outen(`DP5_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_25),
  .pad(`DP5_25),
  .default_value(`default_value)));
ap_DP5_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_25_PULLEN),
  .pullsel(`DP5_25_PULLSEL),
  .pad_pullup(`DP5_25)
));
ap_DP5_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .pullsel(`DP5_25_PULLSEL)
));
ap_DP5_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_25_PULLEN),
  .pullsel(`DP5_25_PULLSEL),
  .pad_pd(`DP5_25)
));
ap_DP5_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_25),
  .pullen(`DP5_25_PULLEN),
  .pullsel(`DP5_25_PULLSEL)
));
ap_DP5_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXCLK_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`RGMII2TXCLK_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXCLK_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`RGMII2TXCLK_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE)
));
ap_DP5_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_26_PINCTRL_0_IE),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_26),
  .pad(`DP5_26),
  .default_value(`default_value)));
ap_DP5_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS3_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`SPI2CS3_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE)
));
ap_DP5_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_26_PINCTRL_0_IE),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_26),
  .pad(`DP5_26),
  .default_value(`default_value)));
ap_DP5_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE)
));
ap_DP5_26_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_26_PINCTRL_0_IE),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_26),
  .pad(`DP5_26),
  .default_value(`default_value)));
ap_DP5_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MCPWM2A_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE)
));
ap_DP5_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_26_PINCTRL_0_IE),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_26),
  .pad(`DP5_26),
  .default_value(`default_value)));
ap_DP5_26_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CLK_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`MIBSPI1CLK_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE)
));
ap_DP5_26_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_26_PINCTRL_0_IE),
  .outen(`DP5_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_26),
  .pad(`DP5_26),
  .default_value(`default_value)));
ap_DP5_26_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP5_26)
));
ap_DP5_26_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_26_OUTFUNC_SEL),
  .gpioouten(`DP5_26_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP5_26_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP5_26),
  .pad_gz(`DP5_26_pad_y)
));
ap_DP5_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_26_PULLEN),
  .pullsel(`DP5_26_PULLSEL),
  .pad_pullup(`DP5_26)
));
ap_DP5_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .pullsel(`DP5_26_PULLSEL)
));
ap_DP5_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_26_PULLEN),
  .pullsel(`DP5_26_PULLSEL),
  .pad_pd(`DP5_26)
));
ap_DP5_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_26),
  .pullen(`DP5_26_PULLEN),
  .pullsel(`DP5_26_PULLSEL)
));
ap_DP5_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD0_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`RGMII2TXD0_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD0_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`RGMII2TXD0_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXCLK_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`FSI1TXCLK_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MCPWM2B_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1PICO_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`MIBSPI1PICO_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_27_OUTFUNC_SEL),
  .gpioouten(`DP5_27_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP5_27_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP5_27),
  .pad_gz(`DP5_27_pad_y)
));
ap_DP5_27_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_27)
));
ap_DP5_27_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE)
));
ap_DP5_27_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_27_PINCTRL_0_IE),
  .outen(`DP5_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_27),
  .pad(`DP5_27),
  .default_value(`default_value)));
ap_DP5_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_27_PULLEN),
  .pullsel(`DP5_27_PULLSEL),
  .pad_pullup(`DP5_27)
));
ap_DP5_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .pullsel(`DP5_27_PULLSEL)
));
ap_DP5_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_27_PULLEN),
  .pullsel(`DP5_27_PULLSEL),
  .pad_pd(`DP5_27)
));
ap_DP5_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_27),
  .pullen(`DP5_27_PULLEN),
  .pullsel(`DP5_27_PULLSEL)
));
ap_DP5_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD1_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`RGMII2TXD1_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD1_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`RGMII2TXD1_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD0_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`FSI1TXD0_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2C_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MCPWM2C_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1POCI_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`MIBSPI1POCI_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_28_OUTFUNC_SEL),
  .gpioouten(`DP5_28_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP5_28_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP5_28),
  .pad_gz(`DP5_28_pad_y)
));
ap_DP5_28_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_28)
));
ap_DP5_28_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE)
));
ap_DP5_28_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_28_PINCTRL_0_IE),
  .outen(`DP5_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_28_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_28),
  .pad(`DP5_28),
  .default_value(`default_value)));
ap_DP5_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_28_PULLEN),
  .pullsel(`DP5_28_PULLSEL),
  .pad_pullup(`DP5_28)
));
ap_DP5_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .pullsel(`DP5_28_PULLSEL)
));
ap_DP5_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_28_PULLEN),
  .pullsel(`DP5_28_PULLSEL),
  .pad_pd(`DP5_28)
));
ap_DP5_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_28),
  .pullen(`DP5_28_PULLEN),
  .pullsel(`DP5_28_PULLSEL)
));
ap_DP5_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD2_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`RGMII2TXD2_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD2_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`RGMII2TXD2_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1TXD1_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`FSI1TXD1_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2D_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MCPWM2D_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_29_OUTFUNC_SEL),
  .gpioouten(`DP5_29_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_29_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_29),
  .pad_gz(`DP5_29_pad_y)
));
ap_DP5_29_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_29)
));
ap_DP5_29_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE)
));
ap_DP5_29_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_29_PINCTRL_0_IE),
  .outen(`DP5_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_29_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_29),
  .pad(`DP5_29),
  .default_value(`default_value)));
ap_DP5_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_29_PULLEN),
  .pullsel(`DP5_29_PULLSEL),
  .pad_pullup(`DP5_29)
));
ap_DP5_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .pullsel(`DP5_29_PULLSEL)
));
ap_DP5_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_29_PULLEN),
  .pullsel(`DP5_29_PULLSEL),
  .pad_pd(`DP5_29)
));
ap_DP5_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_29),
  .pullen(`DP5_29_PULLEN),
  .pullsel(`DP5_29_PULLSEL)
));
ap_DP5_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD3_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`RGMII2TXD3_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXD3_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`RGMII2TXD3_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXCLK_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`FSI1RXCLK_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2E_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MCPWM2E_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_30_OUTFUNC_SEL),
  .gpioouten(`DP5_30_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP5_30_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP5_30),
  .pad_gz(`DP5_30_pad_y)
));
ap_DP5_30_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_30)
));
ap_DP5_30_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE)
));
ap_DP5_30_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_30_PINCTRL_0_IE),
  .outen(`DP5_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_30_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_30),
  .pad(`DP5_30),
  .default_value(`default_value)));
ap_DP5_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_30_PULLEN),
  .pullsel(`DP5_30_PULLSEL),
  .pad_pullup(`DP5_30)
));
ap_DP5_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .pullsel(`DP5_30_PULLSEL)
));
ap_DP5_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_30_PULLEN),
  .pullsel(`DP5_30_PULLSEL),
  .pad_pd(`DP5_30)
));
ap_DP5_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_30),
  .pullen(`DP5_30_PULLEN),
  .pullsel(`DP5_30_PULLSEL)
));
ap_DP5_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXCTL_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`RGMII2TXCTL_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2TXCTL_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`RGMII2TXCTL_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD0_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`FSI1RXD0_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM2F_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MCPWM2F_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CLK_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`SPI9CLK_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP5_31_OUTFUNC_SEL),
  .gpioouten(`DP5_31_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_TX_OE),
  .od(`DP5_31_PINCTRL_0_OD),
  .func_out(`PSI5_2_TX_OUT),
  .pad(`DP5_31),
  .pad_gz(`DP5_31_pad_y)
));
ap_DP5_31_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .pad(`DP5_31)
));
ap_DP5_31_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE)
));
ap_DP5_31_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP5_31_PINCTRL_0_IE),
  .outen(`DP5_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP5_31_INFUNC_EN),
  .in_concat(`input_func_concat_DP5_31),
  .pad(`DP5_31),
  .default_value(`default_value)));
ap_DP5_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP5_31_PULLEN),
  .pullsel(`DP5_31_PULLSEL),
  .pad_pullup(`DP5_31)
));
ap_DP5_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .pullsel(`DP5_31_PULLSEL)
));
ap_DP5_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP5_31_PULLEN),
  .pullsel(`DP5_31_PULLSEL),
  .pad_pd(`DP5_31)
));
ap_DP5_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP5_31),
  .pullen(`DP5_31_PULLEN),
  .pullsel(`DP5_31_PULLSEL)
));
ap_DP6_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXCLK_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`RGMII2RXCLK_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXCLK_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`RGMII2RXCLK_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`FSI1RXD1_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`FSI1RXD1_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3A_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MCPWM3A_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CLK_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`SPI5CLK_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9PICO_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`SPI9PICO_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_0_OUTFUNC_SEL),
  .gpioouten(`DP6_0_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_2_RX_OE),
  .od(`DP6_0_PINCTRL_0_OD),
  .func_out(`PSI5_2_RX_OUT),
  .pad(`DP6_0),
  .pad_gz(`DP6_0_pad_y)
));
ap_DP6_0_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_0)
));
ap_DP6_0_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE)
));
ap_DP6_0_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP6_0_PINCTRL_0_IE),
  .outen(`DP6_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_0),
  .pad(`DP6_0),
  .default_value(`default_value)));
ap_DP6_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_0_PULLEN),
  .pullsel(`DP6_0_PULLSEL),
  .pad_pullup(`DP6_0)
));
ap_DP6_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .pullsel(`DP6_0_PULLSEL)
));
ap_DP6_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_0_PULLEN),
  .pullsel(`DP6_0_PULLSEL),
  .pad_pd(`DP6_0)
));
ap_DP6_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_0),
  .pullen(`DP6_0_PULLEN),
  .pullsel(`DP6_0_PULLSEL)
));
ap_DP6_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD0_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`RGMII2RXD0_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD0_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`RGMII2RXD0_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXCLK_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`FSI2TXCLK_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3B_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`MCPWM3B_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5PICO_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`SPI5PICO_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9POCI_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`SPI9POCI_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_1_OUTFUNC_SEL),
  .gpioouten(`DP6_1_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_TX_OE),
  .od(`DP6_1_PINCTRL_0_OD),
  .func_out(`PSI5_3_TX_OUT),
  .pad(`DP6_1),
  .pad_gz(`DP6_1_pad_y)
));
ap_DP6_1_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_1)
));
ap_DP6_1_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE)
));
ap_DP6_1_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP6_1_PINCTRL_0_IE),
  .outen(`DP6_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_1),
  .pad(`DP6_1),
  .default_value(`default_value)));
ap_DP6_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_1_PULLEN),
  .pullsel(`DP6_1_PULLSEL),
  .pad_pullup(`DP6_1)
));
ap_DP6_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .pullsel(`DP6_1_PULLSEL)
));
ap_DP6_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_1_PULLEN),
  .pullsel(`DP6_1_PULLSEL),
  .pad_pd(`DP6_1)
));
ap_DP6_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_1),
  .pullen(`DP6_1_PULLEN),
  .pullsel(`DP6_1_PULLSEL)
));
ap_DP6_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD1_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`RGMII2RXD1_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD1_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`RGMII2RXD1_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`FSI2TXD0_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3C_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`MCPWM3C_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL0_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5POCI_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`SPI5POCI_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS0_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`SPI9CS0_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_2_OUTFUNC_SEL),
  .gpioouten(`DP6_2_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_3_RX_OE),
  .od(`DP6_2_PINCTRL_0_OD),
  .func_out(`PSI5_3_RX_OUT),
  .pad(`DP6_2),
  .pad_gz(`DP6_2_pad_y)
));
ap_DP6_2_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_2)
));
ap_DP6_2_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE)
));
ap_DP6_2_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP6_2_PINCTRL_0_IE),
  .outen(`DP6_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_2),
  .pad(`DP6_2),
  .default_value(`default_value)));
ap_DP6_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_2_PULLEN),
  .pullsel(`DP6_2_PULLSEL),
  .pad_pullup(`DP6_2)
));
ap_DP6_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .pullsel(`DP6_2_PULLSEL)
));
ap_DP6_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_2_PULLEN),
  .pullsel(`DP6_2_PULLSEL),
  .pad_pd(`DP6_2)
));
ap_DP6_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_2),
  .pullen(`DP6_2_PULLEN),
  .pullsel(`DP6_2_PULLSEL)
));
ap_DP6_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD2_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`RGMII2RXD2_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD2_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`RGMII2RXD2_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2TXD1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`FSI2TXD1_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3D_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`MCPWM3D_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL1_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS0_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`SPI5CS0_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_3_OUTFUNC_SEL),
  .gpioouten(`DP6_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS1_OE),
  .od(`DP6_3_PINCTRL_0_OD),
  .func_out(`SPI9CS1_OUT),
  .pad(`DP6_3),
  .pad_gz(`DP6_3_pad_y)
));
ap_DP6_3_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_3)
));
ap_DP6_3_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE)
));
ap_DP6_3_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_3_PINCTRL_0_IE),
  .outen(`DP6_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_3),
  .pad(`DP6_3),
  .default_value(`default_value)));
ap_DP6_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_3_PULLEN),
  .pullsel(`DP6_3_PULLSEL),
  .pad_pullup(`DP6_3)
));
ap_DP6_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .pullsel(`DP6_3_PULLSEL)
));
ap_DP6_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_3_PULLEN),
  .pullsel(`DP6_3_PULLSEL),
  .pad_pd(`DP6_3)
));
ap_DP6_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_3),
  .pullen(`DP6_3_PULLEN),
  .pullsel(`DP6_3_PULLSEL)
));
ap_DP6_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD3_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`RGMII2RXD3_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXD3_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`RGMII2RXD3_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE)
));
ap_DP6_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_4_PINCTRL_0_IE),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_4),
  .pad(`DP6_4),
  .default_value(`default_value)));
ap_DP6_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC0_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`ADCSOC0_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC0_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`ADCSOC0_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE)
));
ap_DP6_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_4_PINCTRL_0_IE),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_4),
  .pad(`DP6_4),
  .default_value(`default_value)));
ap_DP6_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE)
));
ap_DP6_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_4_PINCTRL_0_IE),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_4),
  .pad(`DP6_4),
  .default_value(`default_value)));
ap_DP6_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3E_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`MCPWM3E_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE)
));
ap_DP6_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_4_PINCTRL_0_IE),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_4),
  .pad(`DP6_4),
  .default_value(`default_value)));
ap_DP6_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL2_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL2_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_4_OUTFUNC_SEL),
  .gpioouten(`DP6_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS2_OE),
  .od(`DP6_4_PINCTRL_0_OD),
  .func_out(`SPI9CS2_OUT),
  .pad(`DP6_4),
  .pad_gz(`DP6_4_pad_y)
));
ap_DP6_4_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_4)
));
ap_DP6_4_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE)
));
ap_DP6_4_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_4_PINCTRL_0_IE),
  .outen(`DP6_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_4),
  .pad(`DP6_4),
  .default_value(`default_value)));
ap_DP6_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_4_PULLEN),
  .pullsel(`DP6_4_PULLSEL),
  .pad_pullup(`DP6_4)
));
ap_DP6_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .pullsel(`DP6_4_PULLSEL)
));
ap_DP6_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_4_PULLEN),
  .pullsel(`DP6_4_PULLSEL),
  .pad_pd(`DP6_4)
));
ap_DP6_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_4),
  .pullen(`DP6_4_PULLEN),
  .pullsel(`DP6_4_PULLSEL)
));
ap_DP6_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXCTL_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`RGMII2RXCTL_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`RGMII2RXCTL_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`RGMII2RXCTL_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE)
));
ap_DP6_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_5_PINCTRL_0_IE),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_5),
  .pad(`DP6_5),
  .default_value(`default_value)));
ap_DP6_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC1_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`ADCSOC1_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADCSOC1_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`ADCSOC1_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE)
));
ap_DP6_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_5_PINCTRL_0_IE),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_5),
  .pad(`DP6_5),
  .default_value(`default_value)));
ap_DP6_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE)
));
ap_DP6_5_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_5_PINCTRL_0_IE),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_5),
  .pad(`DP6_5),
  .default_value(`default_value)));
ap_DP6_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM3F_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`MCPWM3F_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE)
));
ap_DP6_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_5_PINCTRL_0_IE),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_5),
  .pad(`DP6_5),
  .default_value(`default_value)));
ap_DP6_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`ADC5EXTMUXSEL3_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`ADC5EXTMUXSEL3_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_5_OUTFUNC_SEL),
  .gpioouten(`DP6_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS3_OE),
  .od(`DP6_5_PINCTRL_0_OD),
  .func_out(`SPI9CS3_OUT),
  .pad(`DP6_5),
  .pad_gz(`DP6_5_pad_y)
));
ap_DP6_5_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_5)
));
ap_DP6_5_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE)
));
ap_DP6_5_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_5_PINCTRL_0_IE),
  .outen(`DP6_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_5),
  .pad(`DP6_5),
  .default_value(`default_value)));
ap_DP6_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_5_PULLEN),
  .pullsel(`DP6_5_PULLSEL),
  .pad_pullup(`DP6_5)
));
ap_DP6_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .pullsel(`DP6_5_PULLSEL)
));
ap_DP6_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_5_PULLEN),
  .pullsel(`DP6_5_PULLSEL),
  .pad_pd(`DP6_5)
));
ap_DP6_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_5),
  .pullen(`DP6_5_PULLEN),
  .pullsel(`DP6_5_PULLSEL)
));
ap_DP6_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MMC0CLK_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MMC0CLK_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXCLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`FSI2RXCLK_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXCLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`FSI2RXCLK_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MCPWM4A_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1A_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`EPWM1A_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR2_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR2_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_6_OUTFUNC_SEL),
  .gpioouten(`DP6_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`DP6_6_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`DP6_6),
  .pad_gz(`DP6_6_pad_y)
));
ap_DP6_6_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_6)
));
ap_DP6_6_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE)
));
ap_DP6_6_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP6_6_PINCTRL_0_IE),
  .outen(`DP6_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_6),
  .pad(`DP6_6),
  .default_value(`default_value)));
ap_DP6_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_6_PULLEN),
  .pullsel(`DP6_6_PULLSEL),
  .pad_pullup(`DP6_6)
));
ap_DP6_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .pullsel(`DP6_6_PULLSEL)
));
ap_DP6_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_6_PULLEN),
  .pullsel(`DP6_6_PULLSEL),
  .pad_pd(`DP6_6)
));
ap_DP6_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_6),
  .pullen(`DP6_6_PULLEN),
  .pullsel(`DP6_6_PULLSEL)
));
ap_DP6_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CMD_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MMC0CMD_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CMD_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MMC0CMD_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD0_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`FSI2RXD0_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD0_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`FSI2RXD0_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MCPWM4B_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM1B_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`EPWM1B_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR3_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR3_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_8_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_8_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_7_OUTFUNC_SEL),
  .gpioouten(`DP6_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`DP6_7_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`DP6_7),
  .pad_gz(`DP6_7_pad_y)
));
ap_DP6_7_FUNCSEL_8_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_7)
));
ap_DP6_7_FUNCSEL_8_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE)
));
ap_DP6_7_FUNCSEL_8_input_chk : assert property(iomux_input_path(
  .ie(`DP6_7_PINCTRL_0_IE),
  .outen(`DP6_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_7),
  .pad(`DP6_7),
  .default_value(`default_value)));
ap_DP6_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_7_PULLEN),
  .pullsel(`DP6_7_PULLSEL),
  .pad_pullup(`DP6_7)
));
ap_DP6_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .pullsel(`DP6_7_PULLSEL)
));
ap_DP6_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_7_PULLEN),
  .pullsel(`DP6_7_PULLSEL),
  .pad_pd(`DP6_7)
));
ap_DP6_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_7),
  .pullen(`DP6_7_PULLEN),
  .pullsel(`DP6_7_PULLSEL)
));
ap_DP6_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA0_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MMC0DATA0_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA0_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MMC0DATA0_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE)
));
ap_DP6_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_8_PINCTRL_0_IE),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_8),
  .pad(`DP6_8),
  .default_value(`default_value)));
ap_DP6_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD1_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`FSI2RXD1_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`FSI2RXD1_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`FSI2RXD1_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE)
));
ap_DP6_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_8_PINCTRL_0_IE),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_8),
  .pad(`DP6_8),
  .default_value(`default_value)));
ap_DP6_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE)
));
ap_DP6_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_8_PINCTRL_0_IE),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_8),
  .pad(`DP6_8),
  .default_value(`default_value)));
ap_DP6_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4C_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MCPWM4C_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE)
));
ap_DP6_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_8_PINCTRL_0_IE),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_8),
  .pad(`DP6_8),
  .default_value(`default_value)));
ap_DP6_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE)
));
ap_DP6_8_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_8_PINCTRL_0_IE),
  .outen(`DP6_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_8),
  .pad(`DP6_8),
  .default_value(`default_value)));
ap_DP6_8_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2A_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`EPWM2A_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP6_8)
));
ap_DP6_8_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_8_OUTFUNC_SEL),
  .gpioouten(`DP6_8_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR4_OE),
  .od(`DP6_8_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR4_OUT),
  .pad(`DP6_8),
  .pad_gz(`DP6_8_pad_y)
));
ap_DP6_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_8_PULLEN),
  .pullsel(`DP6_8_PULLSEL),
  .pad_pullup(`DP6_8)
));
ap_DP6_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .pullsel(`DP6_8_PULLSEL)
));
ap_DP6_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_8_PULLEN),
  .pullsel(`DP6_8_PULLSEL),
  .pad_pd(`DP6_8)
));
ap_DP6_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_8),
  .pullen(`DP6_8_PULLEN),
  .pullsel(`DP6_8_PULLSEL)
));
ap_DP6_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA1_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MMC0DATA1_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA1_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MMC0DATA1_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE)
));
ap_DP6_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_9_PINCTRL_0_IE),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_9),
  .pad(`DP6_9),
  .default_value(`default_value)));
ap_DP6_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXCLK_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`FSI3TXCLK_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXCLK_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`FSI3TXCLK_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE)
));
ap_DP6_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_9_PINCTRL_0_IE),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_9),
  .pad(`DP6_9),
  .default_value(`default_value)));
ap_DP6_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE)
));
ap_DP6_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_9_PINCTRL_0_IE),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_9),
  .pad(`DP6_9),
  .default_value(`default_value)));
ap_DP6_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4D_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MCPWM4D_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE)
));
ap_DP6_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_9_PINCTRL_0_IE),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_9),
  .pad(`DP6_9),
  .default_value(`default_value)));
ap_DP6_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE)
));
ap_DP6_9_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_9_PINCTRL_0_IE),
  .outen(`DP6_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_9),
  .pad(`DP6_9),
  .default_value(`default_value)));
ap_DP6_9_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM2B_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`EPWM2B_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP6_9)
));
ap_DP6_9_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_9_OUTFUNC_SEL),
  .gpioouten(`DP6_9_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR5_OE),
  .od(`DP6_9_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR5_OUT),
  .pad(`DP6_9),
  .pad_gz(`DP6_9_pad_y)
));
ap_DP6_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_9_PULLEN),
  .pullsel(`DP6_9_PULLSEL),
  .pad_pullup(`DP6_9)
));
ap_DP6_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .pullsel(`DP6_9_PULLSEL)
));
ap_DP6_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_9_PULLEN),
  .pullsel(`DP6_9_PULLSEL),
  .pad_pd(`DP6_9)
));
ap_DP6_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_9),
  .pullen(`DP6_9_PULLEN),
  .pullsel(`DP6_9_PULLSEL)
));
ap_DP6_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA2_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MMC0DATA2_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA2_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MMC0DATA2_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE)
));
ap_DP6_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_10_PINCTRL_0_IE),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_10),
  .pad(`DP6_10),
  .default_value(`default_value)));
ap_DP6_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD0_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`FSI3TXD0_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD0_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`FSI3TXD0_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE)
));
ap_DP6_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_10_PINCTRL_0_IE),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_10),
  .pad(`DP6_10),
  .default_value(`default_value)));
ap_DP6_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE)
));
ap_DP6_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_10_PINCTRL_0_IE),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_10),
  .pad(`DP6_10),
  .default_value(`default_value)));
ap_DP6_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4E_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MCPWM4E_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE)
));
ap_DP6_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_10_PINCTRL_0_IE),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_10),
  .pad(`DP6_10),
  .default_value(`default_value)));
ap_DP6_10_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE)
));
ap_DP6_10_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_10_PINCTRL_0_IE),
  .outen(`DP6_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_10),
  .pad(`DP6_10),
  .default_value(`default_value)));
ap_DP6_10_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3A_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`EPWM3A_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP6_10)
));
ap_DP6_10_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_10_OUTFUNC_SEL),
  .gpioouten(`DP6_10_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR6_OE),
  .od(`DP6_10_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR6_OUT),
  .pad(`DP6_10),
  .pad_gz(`DP6_10_pad_y)
));
ap_DP6_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_10_PULLEN),
  .pullsel(`DP6_10_PULLSEL),
  .pad_pullup(`DP6_10)
));
ap_DP6_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .pullsel(`DP6_10_PULLSEL)
));
ap_DP6_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_10_PULLEN),
  .pullsel(`DP6_10_PULLSEL),
  .pad_pd(`DP6_10)
));
ap_DP6_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_10),
  .pullen(`DP6_10_PULLEN),
  .pullsel(`DP6_10_PULLSEL)
));
ap_DP6_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA3_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MMC0DATA3_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0DATA3_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MMC0DATA3_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE)
));
ap_DP6_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_11_PINCTRL_0_IE),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_11),
  .pad(`DP6_11),
  .default_value(`default_value)));
ap_DP6_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD1_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`FSI3TXD1_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3TXD1_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`FSI3TXD1_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE)
));
ap_DP6_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_11_PINCTRL_0_IE),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_11),
  .pad(`DP6_11),
  .default_value(`default_value)));
ap_DP6_11_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE)
));
ap_DP6_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_11_PINCTRL_0_IE),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_11),
  .pad(`DP6_11),
  .default_value(`default_value)));
ap_DP6_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM4F_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MCPWM4F_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE)
));
ap_DP6_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_11_PINCTRL_0_IE),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_11),
  .pad(`DP6_11),
  .default_value(`default_value)));
ap_DP6_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE)
));
ap_DP6_11_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_11_PINCTRL_0_IE),
  .outen(`DP6_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_11),
  .pad(`DP6_11),
  .default_value(`default_value)));
ap_DP6_11_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM3B_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`EPWM3B_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP6_11)
));
ap_DP6_11_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_11_OUTFUNC_SEL),
  .gpioouten(`DP6_11_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR7_OE),
  .od(`DP6_11_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR7_OUT),
  .pad(`DP6_11),
  .pad_gz(`DP6_11_pad_y)
));
ap_DP6_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_11_PULLEN),
  .pullsel(`DP6_11_PULLSEL),
  .pad_pullup(`DP6_11)
));
ap_DP6_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .pullsel(`DP6_11_PULLSEL)
));
ap_DP6_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_11_PULLEN),
  .pullsel(`DP6_11_PULLSEL),
  .pad_pd(`DP6_11)
));
ap_DP6_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_11),
  .pullen(`DP6_11_PULLEN),
  .pullsel(`DP6_11_PULLSEL)
));
ap_DP6_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CD_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MMC0CD_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0CD_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MMC0CD_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE)
));
ap_DP6_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_12_PINCTRL_0_IE),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_12),
  .pad(`DP6_12),
  .default_value(`default_value)));
ap_DP6_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE)
));
ap_DP6_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_12_PINCTRL_0_IE),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_12),
  .pad(`DP6_12),
  .default_value(`default_value)));
ap_DP6_12_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE)
));
ap_DP6_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_12_PINCTRL_0_IE),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_12),
  .pad(`DP6_12),
  .default_value(`default_value)));
ap_DP6_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5A_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MCPWM5A_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE)
));
ap_DP6_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_12_PINCTRL_0_IE),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_12),
  .pad(`DP6_12),
  .default_value(`default_value)));
ap_DP6_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE)
));
ap_DP6_12_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_12_PINCTRL_0_IE),
  .outen(`DP6_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_12),
  .pad(`DP6_12),
  .default_value(`default_value)));
ap_DP6_12_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP6_12)
));
ap_DP6_12_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_12_OUTFUNC_SEL),
  .gpioouten(`DP6_12_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR8_OE),
  .od(`DP6_12_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR8_OUT),
  .pad(`DP6_12),
  .pad_gz(`DP6_12_pad_y)
));
ap_DP6_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_12_PULLEN),
  .pullsel(`DP6_12_PULLSEL),
  .pad_pullup(`DP6_12)
));
ap_DP6_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .pullsel(`DP6_12_PULLSEL)
));
ap_DP6_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_12_PULLEN),
  .pullsel(`DP6_12_PULLSEL),
  .pad_pd(`DP6_12)
));
ap_DP6_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_12),
  .pullen(`DP6_12_PULLEN),
  .pullsel(`DP6_12_PULLSEL)
));
ap_DP6_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0WP_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MMC0WP_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MMC0WP_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MMC0WP_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE)
));
ap_DP6_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_13_PINCTRL_0_IE),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_13),
  .pad(`DP6_13),
  .default_value(`default_value)));
ap_DP6_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE)
));
ap_DP6_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_13_PINCTRL_0_IE),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_13),
  .pad(`DP6_13),
  .default_value(`default_value)));
ap_DP6_13_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE)
));
ap_DP6_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_13_PINCTRL_0_IE),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_13),
  .pad(`DP6_13),
  .default_value(`default_value)));
ap_DP6_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5B_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`MCPWM5B_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE)
));
ap_DP6_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_13_PINCTRL_0_IE),
  .outen(`DP6_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_13),
  .pad(`DP6_13),
  .default_value(`default_value)));
ap_DP6_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP6_13)
));
ap_DP6_13_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_13_OUTFUNC_SEL),
  .gpioouten(`DP6_13_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR9_OE),
  .od(`DP6_13_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR9_OUT),
  .pad(`DP6_13),
  .pad_gz(`DP6_13_pad_y)
));
ap_DP6_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_13_PULLEN),
  .pullsel(`DP6_13_PULLSEL),
  .pad_pullup(`DP6_13)
));
ap_DP6_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .pullsel(`DP6_13_PULLSEL)
));
ap_DP6_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_13_PULLEN),
  .pullsel(`DP6_13_PULLSEL),
  .pad_pd(`DP6_13)
));
ap_DP6_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_13),
  .pullen(`DP6_13_PULLEN),
  .pullsel(`DP6_13_PULLSEL)
));
ap_DP6_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0TX_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`T1S0TX_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0TX_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`T1S0TX_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE)
));
ap_DP6_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_14_PINCTRL_0_IE),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_14),
  .pad(`DP6_14),
  .default_value(`default_value)));
ap_DP6_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE)
));
ap_DP6_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_14_PINCTRL_0_IE),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_14),
  .pad(`DP6_14),
  .default_value(`default_value)));
ap_DP6_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE)
));
ap_DP6_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_14_PINCTRL_0_IE),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_14),
  .pad(`DP6_14),
  .default_value(`default_value)));
ap_DP6_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5C_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`MCPWM5C_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE)
));
ap_DP6_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_14_PINCTRL_0_IE),
  .outen(`DP6_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_14),
  .pad(`DP6_14),
  .default_value(`default_value)));
ap_DP6_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL0_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL0_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25A_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`EPWM25A_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP6_14)
));
ap_DP6_14_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_14_OUTFUNC_SEL),
  .gpioouten(`DP6_14_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR10_OE),
  .od(`DP6_14_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR10_OUT),
  .pad(`DP6_14),
  .pad_gz(`DP6_14_pad_y)
));
ap_DP6_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_14_PULLEN),
  .pullsel(`DP6_14_PULLSEL),
  .pad_pullup(`DP6_14)
));
ap_DP6_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .pullsel(`DP6_14_PULLSEL)
));
ap_DP6_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_14_PULLEN),
  .pullsel(`DP6_14_PULLSEL),
  .pad_pd(`DP6_14)
));
ap_DP6_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_14),
  .pullen(`DP6_14_PULLEN),
  .pullsel(`DP6_14_PULLSEL)
));
ap_DP6_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0RX_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`T1S0RX_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0RX_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`T1S0RX_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE)
));
ap_DP6_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_15_PINCTRL_0_IE),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_15),
  .pad(`DP6_15),
  .default_value(`default_value)));
ap_DP6_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE)
));
ap_DP6_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_15_PINCTRL_0_IE),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_15),
  .pad(`DP6_15),
  .default_value(`default_value)));
ap_DP6_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE)
));
ap_DP6_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_15_PINCTRL_0_IE),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_15),
  .pad(`DP6_15),
  .default_value(`default_value)));
ap_DP6_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5D_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`MCPWM5D_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE)
));
ap_DP6_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_15_PINCTRL_0_IE),
  .outen(`DP6_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_15),
  .pad(`DP6_15),
  .default_value(`default_value)));
ap_DP6_15_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL1_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL1_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM25B_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`EPWM25B_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP6_15)
));
ap_DP6_15_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_15_OUTFUNC_SEL),
  .gpioouten(`DP6_15_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR11_OE),
  .od(`DP6_15_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR11_OUT),
  .pad(`DP6_15),
  .pad_gz(`DP6_15_pad_y)
));
ap_DP6_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_15_PULLEN),
  .pullsel(`DP6_15_PULLSEL),
  .pad_pullup(`DP6_15)
));
ap_DP6_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .pullsel(`DP6_15_PULLSEL)
));
ap_DP6_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_15_PULLEN),
  .pullsel(`DP6_15_PULLSEL),
  .pad_pd(`DP6_15)
));
ap_DP6_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_15),
  .pullen(`DP6_15_PULLEN),
  .pullsel(`DP6_15_PULLSEL)
));
ap_DP6_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0ED_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`T1S0ED_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`T1S0ED_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`T1S0ED_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE)
));
ap_DP6_16_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_16_PINCTRL_0_IE),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_16),
  .pad(`DP6_16),
  .default_value(`default_value)));
ap_DP6_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE)
));
ap_DP6_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_16_PINCTRL_0_IE),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_16),
  .pad(`DP6_16),
  .default_value(`default_value)));
ap_DP6_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE)
));
ap_DP6_16_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_16_PINCTRL_0_IE),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_16),
  .pad(`DP6_16),
  .default_value(`default_value)));
ap_DP6_16_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5E_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`MCPWM5E_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE)
));
ap_DP6_16_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_16_PINCTRL_0_IE),
  .outen(`DP6_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_16_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_16),
  .pad(`DP6_16),
  .default_value(`default_value)));
ap_DP6_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL2_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL2_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26A_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`EPWM26A_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP6_16)
));
ap_DP6_16_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_16_OUTFUNC_SEL),
  .gpioouten(`DP6_16_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR12_OE),
  .od(`DP6_16_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR12_OUT),
  .pad(`DP6_16),
  .pad_gz(`DP6_16_pad_y)
));
ap_DP6_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_16_PULLEN),
  .pullsel(`DP6_16_PULLSEL),
  .pad_pullup(`DP6_16)
));
ap_DP6_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .pullsel(`DP6_16_PULLSEL)
));
ap_DP6_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_16_PULLEN),
  .pullsel(`DP6_16_PULLSEL),
  .pad_pd(`DP6_16)
));
ap_DP6_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_16),
  .pullen(`DP6_16_PULLEN),
  .pullsel(`DP6_16_PULLSEL)
));
ap_DP6_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1TX_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`T1S1TX_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1TX_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`T1S1TX_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE)
));
ap_DP6_17_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_17_PINCTRL_0_IE),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_17),
  .pad(`DP6_17),
  .default_value(`default_value)));
ap_DP6_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE)
));
ap_DP6_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_17_PINCTRL_0_IE),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_17),
  .pad(`DP6_17),
  .default_value(`default_value)));
ap_DP6_17_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE)
));
ap_DP6_17_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_17_PINCTRL_0_IE),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_17),
  .pad(`DP6_17),
  .default_value(`default_value)));
ap_DP6_17_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM5F_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`MCPWM5F_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE)
));
ap_DP6_17_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_17_PINCTRL_0_IE),
  .outen(`DP6_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_17_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_17),
  .pad(`DP6_17),
  .default_value(`default_value)));
ap_DP6_17_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`ADC4EXTMUXSEL3_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`ADC4EXTMUXSEL3_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM26B_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`EPWM26B_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP6_17)
));
ap_DP6_17_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_17_OUTFUNC_SEL),
  .gpioouten(`DP6_17_GPIO_OUTPUT_ENABLE),
  .oe(`OUTPUTXBAR13_OE),
  .od(`DP6_17_PINCTRL_0_OD),
  .func_out(`OUTPUTXBAR13_OUT),
  .pad(`DP6_17),
  .pad_gz(`DP6_17_pad_y)
));
ap_DP6_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_17_PULLEN),
  .pullsel(`DP6_17_PULLSEL),
  .pad_pullup(`DP6_17)
));
ap_DP6_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .pullsel(`DP6_17_PULLSEL)
));
ap_DP6_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_17_PULLEN),
  .pullsel(`DP6_17_PULLSEL),
  .pad_pd(`DP6_17)
));
ap_DP6_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_17),
  .pullen(`DP6_17_PULLEN),
  .pullsel(`DP6_17_PULLSEL)
));
ap_DP6_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1RX_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`T1S1RX_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1RX_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`T1S1RX_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6A_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MCPWM6A_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT2_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`CLKOUT2_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_18_OUTFUNC_SEL),
  .gpioouten(`DP6_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`DP6_18_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`DP6_18),
  .pad_gz(`DP6_18_pad_y)
));
ap_DP6_18_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_18)
));
ap_DP6_18_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE)
));
ap_DP6_18_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_18_PINCTRL_0_IE),
  .outen(`DP6_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_18_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_18),
  .pad(`DP6_18),
  .default_value(`default_value)));
ap_DP6_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_18_PULLEN),
  .pullsel(`DP6_18_PULLSEL),
  .pad_pullup(`DP6_18)
));
ap_DP6_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .pullsel(`DP6_18_PULLSEL)
));
ap_DP6_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_18_PULLEN),
  .pullsel(`DP6_18_PULLSEL),
  .pad_pd(`DP6_18)
));
ap_DP6_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_18),
  .pullen(`DP6_18_PULLEN),
  .pullsel(`DP6_18_PULLSEL)
));
ap_DP6_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1ED_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`T1S1ED_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`T1S1ED_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`T1S1ED_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`CLKOUT1_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`CLKOUT1_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6B_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MCPWM6B_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CLK_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`SPI3CLK_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_19_OUTFUNC_SEL),
  .gpioouten(`DP6_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`DP6_19_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`DP6_19),
  .pad_gz(`DP6_19_pad_y)
));
ap_DP6_19_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_19)
));
ap_DP6_19_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE)
));
ap_DP6_19_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_19_PINCTRL_0_IE),
  .outen(`DP6_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_19_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_19),
  .pad(`DP6_19),
  .default_value(`default_value)));
ap_DP6_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_19_PULLEN),
  .pullsel(`DP6_19_PULLSEL),
  .pad_pullup(`DP6_19)
));
ap_DP6_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .pullsel(`DP6_19_PULLSEL)
));
ap_DP6_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_19_PULLEN),
  .pullsel(`DP6_19_PULLSEL),
  .pad_pd(`DP6_19)
));
ap_DP6_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_19),
  .pullen(`DP6_19_PULLEN),
  .pullsel(`DP6_19_PULLSEL)
));
ap_DP6_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2TX_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`T1S2TX_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2TX_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`T1S2TX_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CLK_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MSC1CLK_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6C_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MCPWM6C_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3PICO_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`SPI3PICO_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_20_OUTFUNC_SEL),
  .gpioouten(`DP6_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`DP6_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`DP6_20),
  .pad_gz(`DP6_20_pad_y)
));
ap_DP6_20_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_20)
));
ap_DP6_20_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE)
));
ap_DP6_20_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_20_PINCTRL_0_IE),
  .outen(`DP6_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_20_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_20),
  .pad(`DP6_20),
  .default_value(`default_value)));
ap_DP6_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_20_PULLEN),
  .pullsel(`DP6_20_PULLSEL),
  .pad_pullup(`DP6_20)
));
ap_DP6_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .pullsel(`DP6_20_PULLSEL)
));
ap_DP6_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_20_PULLEN),
  .pullsel(`DP6_20_PULLSEL),
  .pad_pd(`DP6_20)
));
ap_DP6_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_20),
  .pullen(`DP6_20_PULLEN),
  .pullsel(`DP6_20_PULLSEL)
));
ap_DP6_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2RX_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`T1S2RX_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2RX_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`T1S2RX_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SI_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MSC1SI_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6D_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MCPWM6D_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3POCI_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`SPI3POCI_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_21_OUTFUNC_SEL),
  .gpioouten(`DP6_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`DP6_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`DP6_21),
  .pad_gz(`DP6_21_pad_y)
));
ap_DP6_21_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_21)
));
ap_DP6_21_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE)
));
ap_DP6_21_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_21_PINCTRL_0_IE),
  .outen(`DP6_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_21_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_21),
  .pad(`DP6_21),
  .default_value(`default_value)));
ap_DP6_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_21_PULLEN),
  .pullsel(`DP6_21_PULLSEL),
  .pad_pullup(`DP6_21)
));
ap_DP6_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .pullsel(`DP6_21_PULLSEL)
));
ap_DP6_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_21_PULLEN),
  .pullsel(`DP6_21_PULLSEL),
  .pad_pd(`DP6_21)
));
ap_DP6_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_21),
  .pullen(`DP6_21_PULLEN),
  .pullsel(`DP6_21_PULLSEL)
));
ap_DP6_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2ED_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`T1S2ED_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`T1S2ED_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`T1S2ED_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1SO_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MSC1SO_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6E_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MCPWM6E_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS0_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`SPI3CS0_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_22_OUTFUNC_SEL),
  .gpioouten(`DP6_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`DP6_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`DP6_22),
  .pad_gz(`DP6_22_pad_y)
));
ap_DP6_22_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_22)
));
ap_DP6_22_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE)
));
ap_DP6_22_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_22_PINCTRL_0_IE),
  .outen(`DP6_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_22_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_22),
  .pad(`DP6_22),
  .default_value(`default_value)));
ap_DP6_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_22_PULLEN),
  .pullsel(`DP6_22_PULLSEL),
  .pad_pullup(`DP6_22)
));
ap_DP6_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .pullsel(`DP6_22_PULLSEL)
));
ap_DP6_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_22_PULLEN),
  .pullsel(`DP6_22_PULLSEL),
  .pad_pd(`DP6_22)
));
ap_DP6_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_22),
  .pullen(`DP6_22_PULLEN),
  .pullsel(`DP6_22_PULLSEL)
));
ap_DP6_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3TX_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`T1S3TX_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3TX_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`T1S3TX_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS0_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MSC1CS0_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM6F_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MCPWM6F_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS1_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`SPI3CS1_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_23_OUTFUNC_SEL),
  .gpioouten(`DP6_23_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`DP6_23_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`DP6_23),
  .pad_gz(`DP6_23_pad_y)
));
ap_DP6_23_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_23)
));
ap_DP6_23_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE)
));
ap_DP6_23_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_23_PINCTRL_0_IE),
  .outen(`DP6_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_23_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_23),
  .pad(`DP6_23),
  .default_value(`default_value)));
ap_DP6_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_23_PULLEN),
  .pullsel(`DP6_23_PULLSEL),
  .pad_pullup(`DP6_23)
));
ap_DP6_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .pullsel(`DP6_23_PULLSEL)
));
ap_DP6_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_23_PULLEN),
  .pullsel(`DP6_23_PULLSEL),
  .pad_pd(`DP6_23)
));
ap_DP6_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_23),
  .pullen(`DP6_23_PULLEN),
  .pullsel(`DP6_23_PULLSEL)
));
ap_DP6_24_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3RX_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`T1S3RX_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3RX_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`T1S3RX_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS1_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MSC1CS1_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7A_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MCPWM7A_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS2_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`SPI3CS2_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_24_OUTFUNC_SEL),
  .gpioouten(`DP6_24_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`DP6_24_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`DP6_24),
  .pad_gz(`DP6_24_pad_y)
));
ap_DP6_24_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_24)
));
ap_DP6_24_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE)
));
ap_DP6_24_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_24_PINCTRL_0_IE),
  .outen(`DP6_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_24_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_24),
  .pad(`DP6_24),
  .default_value(`default_value)));
ap_DP6_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_24_PULLEN),
  .pullsel(`DP6_24_PULLSEL),
  .pad_pullup(`DP6_24)
));
ap_DP6_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .pullsel(`DP6_24_PULLSEL)
));
ap_DP6_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_24_PULLEN),
  .pullsel(`DP6_24_PULLSEL),
  .pad_pd(`DP6_24)
));
ap_DP6_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_24),
  .pullen(`DP6_24_PULLEN),
  .pullsel(`DP6_24_PULLSEL)
));
ap_DP6_25_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3ED_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`T1S3ED_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`T1S3ED_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`T1S3ED_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7B_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MCPWM7B_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS3_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`SPI3CS3_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_7_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_7_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_25_OUTFUNC_SEL),
  .gpioouten(`DP6_25_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`DP6_25_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`DP6_25),
  .pad_gz(`DP6_25_pad_y)
));
ap_DP6_25_FUNCSEL_7_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_25)
));
ap_DP6_25_FUNCSEL_7_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE)
));
ap_DP6_25_FUNCSEL_7_input_chk : assert property(iomux_input_path(
  .ie(`DP6_25_PINCTRL_0_IE),
  .outen(`DP6_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_25_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_25),
  .pad(`DP6_25),
  .default_value(`default_value)));
ap_DP6_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_25_PULLEN),
  .pullsel(`DP6_25_PULLSEL),
  .pad_pullup(`DP6_25)
));
ap_DP6_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .pullsel(`DP6_25_PULLSEL)
));
ap_DP6_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_25_PULLEN),
  .pullsel(`DP6_25_PULLSEL),
  .pad_pd(`DP6_25)
));
ap_DP6_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_25),
  .pullen(`DP6_25_PULLEN),
  .pullsel(`DP6_25_PULLSEL)
));
ap_DP6_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`T1SMDC_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`T1SMDC_OUT),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`T1SMDC_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`T1SMDC_OUT),
  .pad(`DP6_26),
  .pad_gz(`DP6_26_pad_y)
));
ap_DP6_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_26),
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE)
));
ap_DP6_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_26_PINCTRL_0_IE),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_26),
  .pad(`DP6_26),
  .default_value(`default_value)));
ap_DP6_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS2_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`MSC1CS2_OUT),
  .pad(`DP6_26),
  .pad_gz(`DP6_26_pad_y)
));
ap_DP6_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_26),
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE)
));
ap_DP6_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_26_PINCTRL_0_IE),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_26),
  .pad(`DP6_26),
  .default_value(`default_value)));
ap_DP6_26_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL2_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL2_OUT),
  .pad(`DP6_26),
  .pad_gz(`DP6_26_pad_y)
));
ap_DP6_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_26_OUTFUNC_SEL),
  .gpioouten(`DP6_26_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7C_OE),
  .od(`DP6_26_PINCTRL_0_OD),
  .func_out(`MCPWM7C_OUT),
  .pad(`DP6_26),
  .pad_gz(`DP6_26_pad_y)
));
ap_DP6_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_26)
));
ap_DP6_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_26),
  .pullen(`DP6_26_PULLEN),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE)
));
ap_DP6_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_26_PINCTRL_0_IE),
  .outen(`DP6_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_26_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_26),
  .pad(`DP6_26),
  .default_value(`default_value)));
ap_DP6_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_26_PULLEN),
  .pullsel(`DP6_26_PULLSEL),
  .pad_pullup(`DP6_26)
));
ap_DP6_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_26),
  .pullen(`DP6_26_PULLEN),
  .pullsel(`DP6_26_PULLSEL)
));
ap_DP6_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_26_PULLEN),
  .pullsel(`DP6_26_PULLSEL),
  .pad_pd(`DP6_26)
));
ap_DP6_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_26),
  .pullen(`DP6_26_PULLEN),
  .pullsel(`DP6_26_PULLSEL)
));
ap_DP6_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`T1SMDIO_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`T1SMDIO_OUT),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`T1SMDIO_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`T1SMDIO_OUT),
  .pad(`DP6_27),
  .pad_gz(`DP6_27_pad_y)
));
ap_DP6_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_27),
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE)
));
ap_DP6_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP6_27_PINCTRL_0_IE),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_27),
  .pad(`DP6_27),
  .default_value(`default_value)));
ap_DP6_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`MSC1CS3_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`MSC1CS3_OUT),
  .pad(`DP6_27),
  .pad_gz(`DP6_27_pad_y)
));
ap_DP6_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_27),
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE)
));
ap_DP6_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP6_27_PINCTRL_0_IE),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_27),
  .pad(`DP6_27),
  .default_value(`default_value)));
ap_DP6_27_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`ADC6EXTMUXSEL3_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`ADC6EXTMUXSEL3_OUT),
  .pad(`DP6_27),
  .pad_gz(`DP6_27_pad_y)
));
ap_DP6_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP6_27_OUTFUNC_SEL),
  .gpioouten(`DP6_27_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7D_OE),
  .od(`DP6_27_PINCTRL_0_OD),
  .func_out(`MCPWM7D_OUT),
  .pad(`DP6_27),
  .pad_gz(`DP6_27_pad_y)
));
ap_DP6_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .pad(`DP6_27)
));
ap_DP6_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP6_27),
  .pullen(`DP6_27_PULLEN),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE)
));
ap_DP6_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP6_27_PINCTRL_0_IE),
  .outen(`DP6_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP6_27_INFUNC_EN),
  .in_concat(`input_func_concat_DP6_27),
  .pad(`DP6_27),
  .default_value(`default_value)));
ap_DP6_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP6_27_PULLEN),
  .pullsel(`DP6_27_PULLSEL),
  .pad_pullup(`DP6_27)
));
ap_DP6_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP6_27),
  .pullen(`DP6_27_PULLEN),
  .pullsel(`DP6_27_PULLSEL)
));
ap_DP6_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP6_27_PULLEN),
  .pullsel(`DP6_27_PULLSEL),
  .pad_pd(`DP6_27)
));
ap_DP6_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP6_27),
  .pullen(`DP6_27_PULLEN),
  .pullsel(`DP6_27_PULLSEL)
));
ap_DP7_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1A_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1A_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1A_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1A_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0TX_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`LPD_CAN0TX_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0TX_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`LPD_CAN0TX_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CLK_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`MSC0CLK_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE)
));
ap_DP7_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_0_PINCTRL_0_IE),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_0),
  .pad(`DP7_0),
  .default_value(`default_value)));
ap_DP7_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7E_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`MCPWM7E_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE)
));
ap_DP7_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_0_PINCTRL_0_IE),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_0),
  .pad(`DP7_0),
  .default_value(`default_value)));
ap_DP7_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS4_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`SPI2CS4_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE)
));
ap_DP7_0_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_0_PINCTRL_0_IE),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_0),
  .pad(`DP7_0),
  .default_value(`default_value)));
ap_DP7_0_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_0_OUTFUNC_SEL),
  .gpioouten(`DP7_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`DP7_0_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`DP7_0),
  .pad_gz(`DP7_0_pad_y)
));
ap_DP7_0_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_0)
));
ap_DP7_0_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE)
));
ap_DP7_0_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_0_PINCTRL_0_IE),
  .outen(`DP7_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_0_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_0),
  .pad(`DP7_0),
  .default_value(`default_value)));
ap_DP7_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_0_PULLEN),
  .pullsel(`DP7_0_PULLSEL),
  .pad_pullup(`DP7_0)
));
ap_DP7_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .pullsel(`DP7_0_PULLSEL)
));
ap_DP7_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_0_PULLEN),
  .pullsel(`DP7_0_PULLSEL),
  .pad_pd(`DP7_0)
));
ap_DP7_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_0),
  .pullen(`DP7_0_PULLEN),
  .pullsel(`DP7_0_PULLSEL)
));
ap_DP7_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1B_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1B_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1B_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1B_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0RX_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`LPD_CAN0RX_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0RX_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`LPD_CAN0RX_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SI_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`MSC0SI_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE)
));
ap_DP7_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_1_PINCTRL_0_IE),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_1),
  .pad(`DP7_1),
  .default_value(`default_value)));
ap_DP7_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM7F_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`MCPWM7F_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE)
));
ap_DP7_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_1_PINCTRL_0_IE),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_1),
  .pad(`DP7_1),
  .default_value(`default_value)));
ap_DP7_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI2CS5_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`SPI2CS5_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE)
));
ap_DP7_1_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_1_PINCTRL_0_IE),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_1),
  .pad(`DP7_1),
  .default_value(`default_value)));
ap_DP7_1_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_1_OUTFUNC_SEL),
  .gpioouten(`DP7_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`DP7_1_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`DP7_1),
  .pad_gz(`DP7_1_pad_y)
));
ap_DP7_1_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_1)
));
ap_DP7_1_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE)
));
ap_DP7_1_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_1_PINCTRL_0_IE),
  .outen(`DP7_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_1_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_1),
  .pad(`DP7_1),
  .default_value(`default_value)));
ap_DP7_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_1_PULLEN),
  .pullsel(`DP7_1_PULLSEL),
  .pad_pullup(`DP7_1)
));
ap_DP7_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .pullsel(`DP7_1_PULLSEL)
));
ap_DP7_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_1_PULLEN),
  .pullsel(`DP7_1_PULLSEL),
  .pad_pd(`DP7_1)
));
ap_DP7_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_1),
  .pullen(`DP7_1_PULLEN),
  .pullsel(`DP7_1_PULLSEL)
));
ap_DP7_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2A_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2A_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4A_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4A_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0SO_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`MSC0SO_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_2),
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE)
));
ap_DP7_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_2_PINCTRL_0_IE),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_2),
  .pad(`DP7_2),
  .default_value(`default_value)));
ap_DP7_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`MCPWM8A_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_2),
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE)
));
ap_DP7_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_2_PINCTRL_0_IE),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_2),
  .pad(`DP7_2),
  .default_value(`default_value)));
ap_DP7_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21A_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`EPWM21A_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_2_OUTFUNC_SEL),
  .gpioouten(`DP7_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP7_2_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP7_2),
  .pad_gz(`DP7_2_pad_y)
));
ap_DP7_2_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_2)
));
ap_DP7_2_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_2),
  .pullen(`DP7_2_PULLEN),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE)
));
ap_DP7_2_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_2_PINCTRL_0_IE),
  .outen(`DP7_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_2_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_2),
  .pad(`DP7_2),
  .default_value(`default_value)));
ap_DP7_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_2_PULLEN),
  .pullsel(`DP7_2_PULLSEL),
  .pad_pullup(`DP7_2)
));
ap_DP7_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_2),
  .pullen(`DP7_2_PULLEN),
  .pullsel(`DP7_2_PULLSEL)
));
ap_DP7_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_2_PULLEN),
  .pullsel(`DP7_2_PULLSEL),
  .pad_pd(`DP7_2)
));
ap_DP7_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_2),
  .pullen(`DP7_2_PULLEN),
  .pullsel(`DP7_2_PULLSEL)
));
ap_DP7_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2B_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2B_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4B_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4B_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS0_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`MSC0CS0_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_3),
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE)
));
ap_DP7_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_3_PINCTRL_0_IE),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_3),
  .pad(`DP7_3),
  .default_value(`default_value)));
ap_DP7_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`MCPWM8B_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_3),
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE)
));
ap_DP7_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_3_PINCTRL_0_IE),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_3),
  .pad(`DP7_3),
  .default_value(`default_value)));
ap_DP7_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM21B_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`EPWM21B_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_3_OUTFUNC_SEL),
  .gpioouten(`DP7_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP7_3_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP7_3),
  .pad_gz(`DP7_3_pad_y)
));
ap_DP7_3_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_3)
));
ap_DP7_3_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_3),
  .pullen(`DP7_3_PULLEN),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE)
));
ap_DP7_3_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_3_PINCTRL_0_IE),
  .outen(`DP7_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_3_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_3),
  .pad(`DP7_3),
  .default_value(`default_value)));
ap_DP7_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_3_PULLEN),
  .pullsel(`DP7_3_PULLSEL),
  .pad_pullup(`DP7_3)
));
ap_DP7_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_3),
  .pullen(`DP7_3_PULLEN),
  .pullsel(`DP7_3_PULLSEL)
));
ap_DP7_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_3_PULLEN),
  .pullsel(`DP7_3_PULLSEL),
  .pad_pd(`DP7_3)
));
ap_DP7_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_3),
  .pullen(`DP7_3_PULLEN),
  .pullsel(`DP7_3_PULLSEL)
));
ap_DP7_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3A_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3A_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1A_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1A_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS1_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`MSC0CS1_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_4),
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE)
));
ap_DP7_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_4_PINCTRL_0_IE),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_4),
  .pad(`DP7_4),
  .default_value(`default_value)));
ap_DP7_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8C_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`MCPWM8C_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_4),
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE)
));
ap_DP7_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_4_PINCTRL_0_IE),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_4),
  .pad(`DP7_4),
  .default_value(`default_value)));
ap_DP7_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22A_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`EPWM22A_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_4_OUTFUNC_SEL),
  .gpioouten(`DP7_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`DP7_4_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`DP7_4),
  .pad_gz(`DP7_4_pad_y)
));
ap_DP7_4_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_4)
));
ap_DP7_4_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_4),
  .pullen(`DP7_4_PULLEN),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE)
));
ap_DP7_4_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_4_PINCTRL_0_IE),
  .outen(`DP7_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_4_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_4),
  .pad(`DP7_4),
  .default_value(`default_value)));
ap_DP7_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_4_PULLEN),
  .pullsel(`DP7_4_PULLSEL),
  .pad_pullup(`DP7_4)
));
ap_DP7_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_4),
  .pullen(`DP7_4_PULLEN),
  .pullsel(`DP7_4_PULLSEL)
));
ap_DP7_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_4_PULLEN),
  .pullsel(`DP7_4_PULLSEL),
  .pad_pd(`DP7_4)
));
ap_DP7_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_4),
  .pullen(`DP7_4_PULLEN),
  .pullsel(`DP7_4_PULLSEL)
));
ap_DP7_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3B_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3B_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1B_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM1B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM1B_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS2_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`MSC0CS2_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_5),
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE)
));
ap_DP7_5_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_5_PINCTRL_0_IE),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_5),
  .pad(`DP7_5),
  .default_value(`default_value)));
ap_DP7_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8D_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`MCPWM8D_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_5),
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE)
));
ap_DP7_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_5_PINCTRL_0_IE),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_5),
  .pad(`DP7_5),
  .default_value(`default_value)));
ap_DP7_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM22B_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`EPWM22B_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_5_OUTFUNC_SEL),
  .gpioouten(`DP7_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`DP7_5_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`DP7_5),
  .pad_gz(`DP7_5_pad_y)
));
ap_DP7_5_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_5)
));
ap_DP7_5_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_5),
  .pullen(`DP7_5_PULLEN),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE)
));
ap_DP7_5_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_5_PINCTRL_0_IE),
  .outen(`DP7_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_5_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_5),
  .pad(`DP7_5),
  .default_value(`default_value)));
ap_DP7_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_5_PULLEN),
  .pullsel(`DP7_5_PULLSEL),
  .pad_pullup(`DP7_5)
));
ap_DP7_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_5),
  .pullen(`DP7_5_PULLEN),
  .pullsel(`DP7_5_PULLSEL)
));
ap_DP7_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_5_PULLEN),
  .pullsel(`DP7_5_PULLSEL),
  .pad_pd(`DP7_5)
));
ap_DP7_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_5),
  .pullen(`DP7_5_PULLEN),
  .pullsel(`DP7_5_PULLSEL)
));
ap_DP7_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4A_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4A_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2A_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2A_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`MSC0CS3_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`MSC0CS3_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_6),
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE)
));
ap_DP7_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_6_PINCTRL_0_IE),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_6),
  .pad(`DP7_6),
  .default_value(`default_value)));
ap_DP7_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8E_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`MCPWM8E_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_6),
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE)
));
ap_DP7_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_6_PINCTRL_0_IE),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_6),
  .pad(`DP7_6),
  .default_value(`default_value)));
ap_DP7_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23A_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`EPWM23A_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_6_OUTFUNC_SEL),
  .gpioouten(`DP7_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`DP7_6_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`DP7_6),
  .pad_gz(`DP7_6_pad_y)
));
ap_DP7_6_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_6)
));
ap_DP7_6_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_6),
  .pullen(`DP7_6_PULLEN),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE)
));
ap_DP7_6_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_6_PINCTRL_0_IE),
  .outen(`DP7_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_6_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_6),
  .pad(`DP7_6),
  .default_value(`default_value)));
ap_DP7_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_6_PULLEN),
  .pullsel(`DP7_6_PULLSEL),
  .pad_pullup(`DP7_6)
));
ap_DP7_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_6),
  .pullen(`DP7_6_PULLEN),
  .pullsel(`DP7_6_PULLSEL)
));
ap_DP7_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_6_PULLEN),
  .pullsel(`DP7_6_PULLSEL),
  .pad_pd(`DP7_6)
));
ap_DP7_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_6),
  .pullen(`DP7_6_PULLEN),
  .pullsel(`DP7_6_PULLSEL)
));
ap_DP7_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4B_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM4B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM4B_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2B_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_A_PWM2B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`LPD_A_PWM2B_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_TX_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`PSI5_0_TX_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_7),
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE)
));
ap_DP7_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_7_PINCTRL_0_IE),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_7),
  .pad(`DP7_7),
  .default_value(`default_value)));
ap_DP7_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM8F_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`MCPWM8F_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_7),
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE)
));
ap_DP7_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_7_PINCTRL_0_IE),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_7),
  .pad(`DP7_7),
  .default_value(`default_value)));
ap_DP7_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM23B_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`EPWM23B_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_6_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_6_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_7_OUTFUNC_SEL),
  .gpioouten(`DP7_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`DP7_7_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`DP7_7),
  .pad_gz(`DP7_7_pad_y)
));
ap_DP7_7_FUNCSEL_6_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_7)
));
ap_DP7_7_FUNCSEL_6_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_7),
  .pullen(`DP7_7_PULLEN),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE)
));
ap_DP7_7_FUNCSEL_6_input_chk : assert property(iomux_input_path(
  .ie(`DP7_7_PINCTRL_0_IE),
  .outen(`DP7_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_7_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_7),
  .pad(`DP7_7),
  .default_value(`default_value)));
ap_DP7_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_7_PULLEN),
  .pullsel(`DP7_7_PULLSEL),
  .pad_pullup(`DP7_7)
));
ap_DP7_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_7),
  .pullen(`DP7_7_PULLEN),
  .pullsel(`DP7_7_PULLSEL)
));
ap_DP7_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_7_PULLEN),
  .pullsel(`DP7_7_PULLSEL),
  .pad_pd(`DP7_7)
));
ap_DP7_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_7),
  .pullen(`DP7_7_PULLEN),
  .pullsel(`DP7_7_PULLSEL)
));
ap_DP7_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0TX_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`LPD_CAN0TX_OUT),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0TX_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`LPD_CAN0TX_OUT),
  .pad(`DP7_8),
  .pad_gz(`DP7_8_pad_y)
));
ap_DP7_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3A_OUT),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3A_OUT),
  .pad(`DP7_8),
  .pad_gz(`DP7_8_pad_y)
));
ap_DP7_8_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_0_RX_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`PSI5_0_RX_OUT),
  .pad(`DP7_8),
  .pad_gz(`DP7_8_pad_y)
));
ap_DP7_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_8_PULLEN),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_8),
  .pullen(`DP7_8_PULLEN),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE)
));
ap_DP7_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_8_PINCTRL_0_IE),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_8),
  .pad(`DP7_8),
  .default_value(`default_value)));
ap_DP7_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`MCPWM9A_OUT),
  .pad(`DP7_8),
  .pad_gz(`DP7_8_pad_y)
));
ap_DP7_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_8_PULLEN),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_8),
  .pullen(`DP7_8_PULLEN),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE)
));
ap_DP7_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_8_PINCTRL_0_IE),
  .outen(`DP7_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_8_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_8),
  .pad(`DP7_8),
  .default_value(`default_value)));
ap_DP7_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP7_8)
));
ap_DP7_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_8_OUTFUNC_SEL),
  .gpioouten(`DP7_8_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24A_OE),
  .od(`DP7_8_PINCTRL_0_OD),
  .func_out(`EPWM24A_OUT),
  .pad(`DP7_8),
  .pad_gz(`DP7_8_pad_y)
));
ap_DP7_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_8_PULLEN),
  .pullsel(`DP7_8_PULLSEL),
  .pad_pullup(`DP7_8)
));
ap_DP7_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_8),
  .pullen(`DP7_8_PULLEN),
  .pullsel(`DP7_8_PULLSEL)
));
ap_DP7_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_8_PULLEN),
  .pullsel(`DP7_8_PULLSEL),
  .pad_pd(`DP7_8)
));
ap_DP7_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_8),
  .pullen(`DP7_8_PULLEN),
  .pullsel(`DP7_8_PULLSEL)
));
ap_DP7_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0RX_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`LPD_CAN0RX_OUT),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_CAN0RX_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`LPD_CAN0RX_OUT),
  .pad(`DP7_9),
  .pad_gz(`DP7_9_pad_y)
));
ap_DP7_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3B_OUT),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_B_PWM3B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`LPD_B_PWM3B_OUT),
  .pad(`DP7_9),
  .pad_gz(`DP7_9_pad_y)
));
ap_DP7_9_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_TX_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`PSI5_1_TX_OUT),
  .pad(`DP7_9),
  .pad_gz(`DP7_9_pad_y)
));
ap_DP7_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_9_PULLEN),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_9),
  .pullen(`DP7_9_PULLEN),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE)
));
ap_DP7_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_9_PINCTRL_0_IE),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_9),
  .pad(`DP7_9),
  .default_value(`default_value)));
ap_DP7_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`MCPWM9B_OUT),
  .pad(`DP7_9),
  .pad_gz(`DP7_9_pad_y)
));
ap_DP7_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_9_PULLEN),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_9),
  .pullen(`DP7_9_PULLEN),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE)
));
ap_DP7_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_9_PINCTRL_0_IE),
  .outen(`DP7_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_9_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_9),
  .pad(`DP7_9),
  .default_value(`default_value)));
ap_DP7_9_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP7_9)
));
ap_DP7_9_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_9_OUTFUNC_SEL),
  .gpioouten(`DP7_9_GPIO_OUTPUT_ENABLE),
  .oe(`EPWM24B_OE),
  .od(`DP7_9_PINCTRL_0_OD),
  .func_out(`EPWM24B_OUT),
  .pad(`DP7_9),
  .pad_gz(`DP7_9_pad_y)
));
ap_DP7_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_9_PULLEN),
  .pullsel(`DP7_9_PULLSEL),
  .pad_pullup(`DP7_9)
));
ap_DP7_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_9),
  .pullen(`DP7_9_PULLEN),
  .pullsel(`DP7_9_PULLSEL)
));
ap_DP7_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_9_PULLEN),
  .pullsel(`DP7_9_PULLSEL),
  .pad_pd(`DP7_9)
));
ap_DP7_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_9),
  .pullen(`DP7_9_PULLEN),
  .pullsel(`DP7_9_PULLSEL)
));
ap_DP7_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_10)
));
ap_DP7_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_10),
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE)
));
ap_DP7_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_10_PINCTRL_0_IE),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_10),
  .pad(`DP7_10),
  .default_value(`default_value)));
ap_DP7_10_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_10_OUTFUNC_SEL),
  .gpioouten(`DP7_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP7_10_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP7_10)
));
ap_DP7_10_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_10_OUTFUNC_SEL),
  .gpioouten(`DP7_10_GPIO_OUTPUT_ENABLE),
  .oe(`PSI5_1_RX_OE),
  .od(`DP7_10_PINCTRL_0_OD),
  .func_out(`PSI5_1_RX_OUT),
  .pad(`DP7_10),
  .pad_gz(`DP7_10_pad_y)
));
ap_DP7_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_10)
));
ap_DP7_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_10),
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE)
));
ap_DP7_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`DP7_10_PINCTRL_0_IE),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_10),
  .pad(`DP7_10),
  .default_value(`default_value)));
ap_DP7_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_10_OUTFUNC_SEL),
  .gpioouten(`DP7_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP7_10_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP7_10)
));
ap_DP7_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_10_OUTFUNC_SEL),
  .gpioouten(`DP7_10_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9C_OE),
  .od(`DP7_10_PINCTRL_0_OD),
  .func_out(`MCPWM9C_OUT),
  .pad(`DP7_10),
  .pad_gz(`DP7_10_pad_y)
));
ap_DP7_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_10)
));
ap_DP7_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_10),
  .pullen(`DP7_10_PULLEN),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE)
));
ap_DP7_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_10_PINCTRL_0_IE),
  .outen(`DP7_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_10_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_10),
  .pad(`DP7_10),
  .default_value(`default_value)));
ap_DP7_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_10_PULLEN),
  .pullsel(`DP7_10_PULLSEL),
  .pad_pullup(`DP7_10)
));
ap_DP7_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_10),
  .pullen(`DP7_10_PULLEN),
  .pullsel(`DP7_10_PULLSEL)
));
ap_DP7_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_10_PULLEN),
  .pullsel(`DP7_10_PULLSEL),
  .pad_pd(`DP7_10)
));
ap_DP7_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_10),
  .pullen(`DP7_10_PULLEN),
  .pullsel(`DP7_10_PULLSEL)
));
ap_DP7_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE)
));
ap_DP7_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_11_PINCTRL_0_IE),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_11),
  .pad(`DP7_11),
  .default_value(`default_value)));
ap_DP7_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`DP7_11),
  .pad_gz(`DP7_11_pad_y)
));
ap_DP7_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE)
));
ap_DP7_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP7_11_PINCTRL_0_IE),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_11),
  .pad(`DP7_11),
  .default_value(`default_value)));
ap_DP7_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9D_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`MCPWM9D_OUT),
  .pad(`DP7_11),
  .pad_gz(`DP7_11_pad_y)
));
ap_DP7_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE)
));
ap_DP7_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_11_PINCTRL_0_IE),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_11),
  .pad(`DP7_11),
  .default_value(`default_value)));
ap_DP7_11_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_11_OUTFUNC_SEL),
  .gpioouten(`DP7_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`DP7_11_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`DP7_11),
  .pad_gz(`DP7_11_pad_y)
));
ap_DP7_11_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_11)
));
ap_DP7_11_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE)
));
ap_DP7_11_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_11_PINCTRL_0_IE),
  .outen(`DP7_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_11_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_11),
  .pad(`DP7_11),
  .default_value(`default_value)));
ap_DP7_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_11_PULLEN),
  .pullsel(`DP7_11_PULLSEL),
  .pad_pullup(`DP7_11)
));
ap_DP7_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .pullsel(`DP7_11_PULLSEL)
));
ap_DP7_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_11_PULLEN),
  .pullsel(`DP7_11_PULLSEL),
  .pad_pd(`DP7_11)
));
ap_DP7_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_11),
  .pullen(`DP7_11_PULLEN),
  .pullsel(`DP7_11_PULLSEL)
));
ap_DP7_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE)
));
ap_DP7_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_12_PINCTRL_0_IE),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_12),
  .pad(`DP7_12),
  .default_value(`default_value)));
ap_DP7_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`DP7_12),
  .pad_gz(`DP7_12_pad_y)
));
ap_DP7_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE)
));
ap_DP7_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP7_12_PINCTRL_0_IE),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_12),
  .pad(`DP7_12),
  .default_value(`default_value)));
ap_DP7_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9E_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`MCPWM9E_OUT),
  .pad(`DP7_12),
  .pad_gz(`DP7_12_pad_y)
));
ap_DP7_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE)
));
ap_DP7_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_12_PINCTRL_0_IE),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_12),
  .pad(`DP7_12),
  .default_value(`default_value)));
ap_DP7_12_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_12_OUTFUNC_SEL),
  .gpioouten(`DP7_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`DP7_12_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`DP7_12),
  .pad_gz(`DP7_12_pad_y)
));
ap_DP7_12_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_12)
));
ap_DP7_12_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE)
));
ap_DP7_12_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_12_PINCTRL_0_IE),
  .outen(`DP7_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_12_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_12),
  .pad(`DP7_12),
  .default_value(`default_value)));
ap_DP7_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_12_PULLEN),
  .pullsel(`DP7_12_PULLSEL),
  .pad_pullup(`DP7_12)
));
ap_DP7_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .pullsel(`DP7_12_PULLSEL)
));
ap_DP7_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_12_PULLEN),
  .pullsel(`DP7_12_PULLSEL),
  .pad_pd(`DP7_12)
));
ap_DP7_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_12),
  .pullen(`DP7_12_PULLEN),
  .pullsel(`DP7_12_PULLSEL)
));
ap_DP7_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE)
));
ap_DP7_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_13_PINCTRL_0_IE),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_13),
  .pad(`DP7_13),
  .default_value(`default_value)));
ap_DP7_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXCLK_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`FSI3RXCLK_OUT),
  .pad(`DP7_13),
  .pad_gz(`DP7_13_pad_y)
));
ap_DP7_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE)
));
ap_DP7_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP7_13_PINCTRL_0_IE),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_13),
  .pad(`DP7_13),
  .default_value(`default_value)));
ap_DP7_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM9F_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`MCPWM9F_OUT),
  .pad(`DP7_13),
  .pad_gz(`DP7_13_pad_y)
));
ap_DP7_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE)
));
ap_DP7_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_13_PINCTRL_0_IE),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_13),
  .pad(`DP7_13),
  .default_value(`default_value)));
ap_DP7_13_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_13_OUTFUNC_SEL),
  .gpioouten(`DP7_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`DP7_13_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`DP7_13),
  .pad_gz(`DP7_13_pad_y)
));
ap_DP7_13_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_13)
));
ap_DP7_13_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE)
));
ap_DP7_13_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_13_PINCTRL_0_IE),
  .outen(`DP7_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_13_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_13),
  .pad(`DP7_13),
  .default_value(`default_value)));
ap_DP7_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_13_PULLEN),
  .pullsel(`DP7_13_PULLSEL),
  .pad_pullup(`DP7_13)
));
ap_DP7_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .pullsel(`DP7_13_PULLSEL)
));
ap_DP7_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_13_PULLEN),
  .pullsel(`DP7_13_PULLSEL),
  .pad_pd(`DP7_13)
));
ap_DP7_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_13),
  .pullen(`DP7_13_PULLEN),
  .pullsel(`DP7_13_PULLSEL)
));
ap_DP7_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE)
));
ap_DP7_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_14_PINCTRL_0_IE),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_14),
  .pad(`DP7_14),
  .default_value(`default_value)));
ap_DP7_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD0_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`FSI3RXD0_OUT),
  .pad(`DP7_14),
  .pad_gz(`DP7_14_pad_y)
));
ap_DP7_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE)
));
ap_DP7_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP7_14_PINCTRL_0_IE),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_14),
  .pad(`DP7_14),
  .default_value(`default_value)));
ap_DP7_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10A_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`MCPWM10A_OUT),
  .pad(`DP7_14),
  .pad_gz(`DP7_14_pad_y)
));
ap_DP7_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE)
));
ap_DP7_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_14_PINCTRL_0_IE),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_14),
  .pad(`DP7_14),
  .default_value(`default_value)));
ap_DP7_14_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_14_OUTFUNC_SEL),
  .gpioouten(`DP7_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`DP7_14_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`DP7_14),
  .pad_gz(`DP7_14_pad_y)
));
ap_DP7_14_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_14)
));
ap_DP7_14_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE)
));
ap_DP7_14_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`DP7_14_PINCTRL_0_IE),
  .outen(`DP7_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_14_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_14),
  .pad(`DP7_14),
  .default_value(`default_value)));
ap_DP7_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_14_PULLEN),
  .pullsel(`DP7_14_PULLSEL),
  .pad_pullup(`DP7_14)
));
ap_DP7_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .pullsel(`DP7_14_PULLSEL)
));
ap_DP7_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_14_PULLEN),
  .pullsel(`DP7_14_PULLSEL),
  .pad_pd(`DP7_14)
));
ap_DP7_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_14),
  .pullen(`DP7_14_PULLEN),
  .pullsel(`DP7_14_PULLSEL)
));
ap_DP7_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_15)
));
ap_DP7_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_15),
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE)
));
ap_DP7_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`DP7_15_PINCTRL_0_IE),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_15),
  .pad(`DP7_15),
  .default_value(`default_value)));
ap_DP7_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_15_OUTFUNC_SEL),
  .gpioouten(`DP7_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP7_15_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP7_15)
));
ap_DP7_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_15_OUTFUNC_SEL),
  .gpioouten(`DP7_15_GPIO_OUTPUT_ENABLE),
  .oe(`FSI3RXD1_OE),
  .od(`DP7_15_PINCTRL_0_OD),
  .func_out(`FSI3RXD1_OUT),
  .pad(`DP7_15),
  .pad_gz(`DP7_15_pad_y)
));
ap_DP7_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_15)
));
ap_DP7_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_15),
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE)
));
ap_DP7_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`DP7_15_PINCTRL_0_IE),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_15),
  .pad(`DP7_15),
  .default_value(`default_value)));
ap_DP7_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`DP7_15_OUTFUNC_SEL),
  .gpioouten(`DP7_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP7_15_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP7_15)
));
ap_DP7_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`DP7_15_OUTFUNC_SEL),
  .gpioouten(`DP7_15_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10B_OE),
  .od(`DP7_15_PINCTRL_0_OD),
  .func_out(`MCPWM10B_OUT),
  .pad(`DP7_15),
  .pad_gz(`DP7_15_pad_y)
));
ap_DP7_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .pad(`DP7_15)
));
ap_DP7_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`DP7_15),
  .pullen(`DP7_15_PULLEN),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE)
));
ap_DP7_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`DP7_15_PINCTRL_0_IE),
  .outen(`DP7_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`DP7_15_INFUNC_EN),
  .in_concat(`input_func_concat_DP7_15),
  .pad(`DP7_15),
  .default_value(`default_value)));
ap_DP7_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`DP7_15_PULLEN),
  .pullsel(`DP7_15_PULLSEL),
  .pad_pullup(`DP7_15)
));
ap_DP7_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`DP7_15),
  .pullen(`DP7_15_PULLEN),
  .pullsel(`DP7_15_PULLSEL)
));
ap_DP7_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`DP7_15_PULLEN),
  .pullsel(`DP7_15_PULLSEL),
  .pad_pd(`DP7_15)
));
ap_DP7_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`DP7_15),
  .pullen(`DP7_15_PULLEN),
  .pullsel(`DP7_15_PULLSEL)
));
ap_MP2_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE)
));
ap_MP2_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_0_PINCTRL_0_IE),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_0),
  .pad(`MP2_0),
  .default_value(`default_value)));
ap_MP2_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0TX_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`CAN0TX_OUT),
  .pad(`MP2_0),
  .pad_gz(`MP2_0_pad_y)
));
ap_MP2_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE)
));
ap_MP2_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_0_PINCTRL_0_IE),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_0),
  .pad(`MP2_0),
  .default_value(`default_value)));
ap_MP2_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`MP2_0),
  .pad_gz(`MP2_0_pad_y)
));
ap_MP2_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE)
));
ap_MP2_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_0_PINCTRL_0_IE),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_0),
  .pad(`MP2_0),
  .default_value(`default_value)));
ap_MP2_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10C_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`MCPWM10C_OUT),
  .pad(`MP2_0),
  .pad_gz(`MP2_0_pad_y)
));
ap_MP2_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE)
));
ap_MP2_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_0_PINCTRL_0_IE),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_0),
  .pad(`MP2_0),
  .default_value(`default_value)));
ap_MP2_0_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_0_OUTFUNC_SEL),
  .gpioouten(`MP2_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP2_0_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP2_0),
  .pad_gz(`MP2_0_pad_y)
));
ap_MP2_0_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_0)
));
ap_MP2_0_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE)
));
ap_MP2_0_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_0_PINCTRL_0_IE),
  .outen(`MP2_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_0),
  .pad(`MP2_0),
  .default_value(`default_value)));
ap_MP2_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_0_PULLEN),
  .pullsel(`MP2_0_PULLSEL),
  .pad_pullup(`MP2_0)
));
ap_MP2_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .pullsel(`MP2_0_PULLSEL)
));
ap_MP2_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_0_PULLEN),
  .pullsel(`MP2_0_PULLSEL),
  .pad_pd(`MP2_0)
));
ap_MP2_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_0),
  .pullen(`MP2_0_PULLEN),
  .pullsel(`MP2_0_PULLSEL)
));
ap_MP2_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE)
));
ap_MP2_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_1_PINCTRL_0_IE),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_1),
  .pad(`MP2_1),
  .default_value(`default_value)));
ap_MP2_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN0RX_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`CAN0RX_OUT),
  .pad(`MP2_1),
  .pad_gz(`MP2_1_pad_y)
));
ap_MP2_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE)
));
ap_MP2_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_1_PINCTRL_0_IE),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_1),
  .pad(`MP2_1),
  .default_value(`default_value)));
ap_MP2_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`MP2_1),
  .pad_gz(`MP2_1_pad_y)
));
ap_MP2_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE)
));
ap_MP2_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_1_PINCTRL_0_IE),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_1),
  .pad(`MP2_1),
  .default_value(`default_value)));
ap_MP2_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10D_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`MCPWM10D_OUT),
  .pad(`MP2_1),
  .pad_gz(`MP2_1_pad_y)
));
ap_MP2_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE)
));
ap_MP2_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_1_PINCTRL_0_IE),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_1),
  .pad(`MP2_1),
  .default_value(`default_value)));
ap_MP2_1_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_1_OUTFUNC_SEL),
  .gpioouten(`MP2_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP2_1_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP2_1),
  .pad_gz(`MP2_1_pad_y)
));
ap_MP2_1_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_1)
));
ap_MP2_1_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE)
));
ap_MP2_1_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_1_PINCTRL_0_IE),
  .outen(`MP2_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_1),
  .pad(`MP2_1),
  .default_value(`default_value)));
ap_MP2_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_1_PULLEN),
  .pullsel(`MP2_1_PULLSEL),
  .pad_pullup(`MP2_1)
));
ap_MP2_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .pullsel(`MP2_1_PULLSEL)
));
ap_MP2_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_1_PULLEN),
  .pullsel(`MP2_1_PULLSEL),
  .pad_pd(`MP2_1)
));
ap_MP2_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_1),
  .pullen(`MP2_1_PULLEN),
  .pullsel(`MP2_1_PULLSEL)
));
ap_MP2_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE)
));
ap_MP2_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_2_PINCTRL_0_IE),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_2),
  .pad(`MP2_2),
  .default_value(`default_value)));
ap_MP2_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1TX_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`CAN1TX_OUT),
  .pad(`MP2_2),
  .pad_gz(`MP2_2_pad_y)
));
ap_MP2_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE)
));
ap_MP2_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_2_PINCTRL_0_IE),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_2),
  .pad(`MP2_2),
  .default_value(`default_value)));
ap_MP2_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`MP2_2),
  .pad_gz(`MP2_2_pad_y)
));
ap_MP2_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE)
));
ap_MP2_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_2_PINCTRL_0_IE),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_2),
  .pad(`MP2_2),
  .default_value(`default_value)));
ap_MP2_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10E_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`MCPWM10E_OUT),
  .pad(`MP2_2),
  .pad_gz(`MP2_2_pad_y)
));
ap_MP2_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE)
));
ap_MP2_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_2_PINCTRL_0_IE),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_2),
  .pad(`MP2_2),
  .default_value(`default_value)));
ap_MP2_2_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_2_OUTFUNC_SEL),
  .gpioouten(`MP2_2_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP2_2_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP2_2),
  .pad_gz(`MP2_2_pad_y)
));
ap_MP2_2_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_2)
));
ap_MP2_2_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE)
));
ap_MP2_2_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_2_PINCTRL_0_IE),
  .outen(`MP2_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_2),
  .pad(`MP2_2),
  .default_value(`default_value)));
ap_MP2_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_2_PULLEN),
  .pullsel(`MP2_2_PULLSEL),
  .pad_pullup(`MP2_2)
));
ap_MP2_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .pullsel(`MP2_2_PULLSEL)
));
ap_MP2_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_2_PULLEN),
  .pullsel(`MP2_2_PULLSEL),
  .pad_pd(`MP2_2)
));
ap_MP2_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_2),
  .pullen(`MP2_2_PULLEN),
  .pullsel(`MP2_2_PULLSEL)
));
ap_MP2_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE)
));
ap_MP2_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_3_PINCTRL_0_IE),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_3),
  .pad(`MP2_3),
  .default_value(`default_value)));
ap_MP2_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN1RX_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`CAN1RX_OUT),
  .pad(`MP2_3),
  .pad_gz(`MP2_3_pad_y)
));
ap_MP2_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE)
));
ap_MP2_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_3_PINCTRL_0_IE),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_3),
  .pad(`MP2_3),
  .default_value(`default_value)));
ap_MP2_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`MP2_3),
  .pad_gz(`MP2_3_pad_y)
));
ap_MP2_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE)
));
ap_MP2_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_3_PINCTRL_0_IE),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_3),
  .pad(`MP2_3),
  .default_value(`default_value)));
ap_MP2_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`MCPWM10F_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`MCPWM10F_OUT),
  .pad(`MP2_3),
  .pad_gz(`MP2_3_pad_y)
));
ap_MP2_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE)
));
ap_MP2_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_3_PINCTRL_0_IE),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_3),
  .pad(`MP2_3),
  .default_value(`default_value)));
ap_MP2_3_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_3_OUTFUNC_SEL),
  .gpioouten(`MP2_3_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP2_3_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP2_3),
  .pad_gz(`MP2_3_pad_y)
));
ap_MP2_3_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_3)
));
ap_MP2_3_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE)
));
ap_MP2_3_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_3_PINCTRL_0_IE),
  .outen(`MP2_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_3),
  .pad(`MP2_3),
  .default_value(`default_value)));
ap_MP2_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_3_PULLEN),
  .pullsel(`MP2_3_PULLSEL),
  .pad_pullup(`MP2_3)
));
ap_MP2_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .pullsel(`MP2_3_PULLSEL)
));
ap_MP2_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_3_PULLEN),
  .pullsel(`MP2_3_PULLSEL),
  .pad_pd(`MP2_3)
));
ap_MP2_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_3),
  .pullen(`MP2_3_PULLEN),
  .pullsel(`MP2_3_PULLSEL)
));
ap_MP2_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE)
));
ap_MP2_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_4_PINCTRL_0_IE),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_4),
  .pad(`MP2_4),
  .default_value(`default_value)));
ap_MP2_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2TX_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`CAN2TX_OUT),
  .pad(`MP2_4),
  .pad_gz(`MP2_4_pad_y)
));
ap_MP2_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE)
));
ap_MP2_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_4_PINCTRL_0_IE),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_4),
  .pad(`MP2_4),
  .default_value(`default_value)));
ap_MP2_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`MP2_4),
  .pad_gz(`MP2_4_pad_y)
));
ap_MP2_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE)
));
ap_MP2_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_4_PINCTRL_0_IE),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_4),
  .pad(`MP2_4),
  .default_value(`default_value)));
ap_MP2_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`MP2_4),
  .pad_gz(`MP2_4_pad_y)
));
ap_MP2_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE)
));
ap_MP2_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_4_PINCTRL_0_IE),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_4),
  .pad(`MP2_4),
  .default_value(`default_value)));
ap_MP2_4_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_4_OUTFUNC_SEL),
  .gpioouten(`MP2_4_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_N_OE),
  .od(`MP2_4_PINCTRL_0_OD),
  .func_out(`RDC0PWM_N_OUT),
  .pad(`MP2_4),
  .pad_gz(`MP2_4_pad_y)
));
ap_MP2_4_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_4)
));
ap_MP2_4_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE)
));
ap_MP2_4_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_4_PINCTRL_0_IE),
  .outen(`MP2_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_4),
  .pad(`MP2_4),
  .default_value(`default_value)));
ap_MP2_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_4_PULLEN),
  .pullsel(`MP2_4_PULLSEL),
  .pad_pullup(`MP2_4)
));
ap_MP2_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .pullsel(`MP2_4_PULLSEL)
));
ap_MP2_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_4_PULLEN),
  .pullsel(`MP2_4_PULLSEL),
  .pad_pd(`MP2_4)
));
ap_MP2_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_4),
  .pullen(`MP2_4_PULLEN),
  .pullsel(`MP2_4_PULLSEL)
));
ap_MP2_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE)
));
ap_MP2_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_5_PINCTRL_0_IE),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_5),
  .pad(`MP2_5),
  .default_value(`default_value)));
ap_MP2_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN2RX_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`CAN2RX_OUT),
  .pad(`MP2_5),
  .pad_gz(`MP2_5_pad_y)
));
ap_MP2_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE)
));
ap_MP2_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_5_PINCTRL_0_IE),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_5),
  .pad(`MP2_5),
  .default_value(`default_value)));
ap_MP2_5_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`MP2_5),
  .pad_gz(`MP2_5_pad_y)
));
ap_MP2_5_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE)
));
ap_MP2_5_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_5_PINCTRL_0_IE),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_5),
  .pad(`MP2_5),
  .default_value(`default_value)));
ap_MP2_5_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`MP2_5),
  .pad_gz(`MP2_5_pad_y)
));
ap_MP2_5_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE)
));
ap_MP2_5_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_5_PINCTRL_0_IE),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_5),
  .pad(`MP2_5),
  .default_value(`default_value)));
ap_MP2_5_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_5_OUTFUNC_SEL),
  .gpioouten(`MP2_5_GPIO_OUTPUT_ENABLE),
  .oe(`RDC0PWM_P_OE),
  .od(`MP2_5_PINCTRL_0_OD),
  .func_out(`RDC0PWM_P_OUT),
  .pad(`MP2_5),
  .pad_gz(`MP2_5_pad_y)
));
ap_MP2_5_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_5)
));
ap_MP2_5_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE)
));
ap_MP2_5_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_5_PINCTRL_0_IE),
  .outen(`MP2_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_5),
  .pad(`MP2_5),
  .default_value(`default_value)));
ap_MP2_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_5_PULLEN),
  .pullsel(`MP2_5_PULLSEL),
  .pad_pullup(`MP2_5)
));
ap_MP2_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .pullsel(`MP2_5_PULLSEL)
));
ap_MP2_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_5_PULLEN),
  .pullsel(`MP2_5_PULLSEL),
  .pad_pd(`MP2_5)
));
ap_MP2_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_5),
  .pullen(`MP2_5_PULLEN),
  .pullsel(`MP2_5_PULLSEL)
));
ap_MP2_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE)
));
ap_MP2_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_6_PINCTRL_0_IE),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_6),
  .pad(`MP2_6),
  .default_value(`default_value)));
ap_MP2_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3TX_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`CAN3TX_OUT),
  .pad(`MP2_6),
  .pad_gz(`MP2_6_pad_y)
));
ap_MP2_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE)
));
ap_MP2_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_6_PINCTRL_0_IE),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_6),
  .pad(`MP2_6),
  .default_value(`default_value)));
ap_MP2_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`MP2_6),
  .pad_gz(`MP2_6_pad_y)
));
ap_MP2_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE)
));
ap_MP2_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_6_PINCTRL_0_IE),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_6),
  .pad(`MP2_6),
  .default_value(`default_value)));
ap_MP2_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`MP2_6),
  .pad_gz(`MP2_6_pad_y)
));
ap_MP2_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE)
));
ap_MP2_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_6_PINCTRL_0_IE),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_6),
  .pad(`MP2_6),
  .default_value(`default_value)));
ap_MP2_6_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_6_OUTFUNC_SEL),
  .gpioouten(`MP2_6_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_N_OE),
  .od(`MP2_6_PINCTRL_0_OD),
  .func_out(`RDC1PWM_N_OUT),
  .pad(`MP2_6),
  .pad_gz(`MP2_6_pad_y)
));
ap_MP2_6_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_6)
));
ap_MP2_6_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE)
));
ap_MP2_6_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_6_PINCTRL_0_IE),
  .outen(`MP2_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_6),
  .pad(`MP2_6),
  .default_value(`default_value)));
ap_MP2_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_6_PULLEN),
  .pullsel(`MP2_6_PULLSEL),
  .pad_pullup(`MP2_6)
));
ap_MP2_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .pullsel(`MP2_6_PULLSEL)
));
ap_MP2_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_6_PULLEN),
  .pullsel(`MP2_6_PULLSEL),
  .pad_pd(`MP2_6)
));
ap_MP2_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_6),
  .pullen(`MP2_6_PULLEN),
  .pullsel(`MP2_6_PULLSEL)
));
ap_MP2_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE)
));
ap_MP2_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_7_PINCTRL_0_IE),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_7),
  .pad(`MP2_7),
  .default_value(`default_value)));
ap_MP2_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN3RX_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`CAN3RX_OUT),
  .pad(`MP2_7),
  .pad_gz(`MP2_7_pad_y)
));
ap_MP2_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE)
));
ap_MP2_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_7_PINCTRL_0_IE),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_7),
  .pad(`MP2_7),
  .default_value(`default_value)));
ap_MP2_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`MP2_7),
  .pad_gz(`MP2_7_pad_y)
));
ap_MP2_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE)
));
ap_MP2_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_7_PINCTRL_0_IE),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_7),
  .pad(`MP2_7),
  .default_value(`default_value)));
ap_MP2_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`MP2_7),
  .pad_gz(`MP2_7_pad_y)
));
ap_MP2_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE)
));
ap_MP2_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_7_PINCTRL_0_IE),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_7),
  .pad(`MP2_7),
  .default_value(`default_value)));
ap_MP2_7_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_7_OUTFUNC_SEL),
  .gpioouten(`MP2_7_GPIO_OUTPUT_ENABLE),
  .oe(`RDC1PWM_P_OE),
  .od(`MP2_7_PINCTRL_0_OD),
  .func_out(`RDC1PWM_P_OUT),
  .pad(`MP2_7),
  .pad_gz(`MP2_7_pad_y)
));
ap_MP2_7_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_7)
));
ap_MP2_7_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE)
));
ap_MP2_7_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP2_7_PINCTRL_0_IE),
  .outen(`MP2_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_7),
  .pad(`MP2_7),
  .default_value(`default_value)));
ap_MP2_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_7_PULLEN),
  .pullsel(`MP2_7_PULLSEL),
  .pad_pullup(`MP2_7)
));
ap_MP2_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .pullsel(`MP2_7_PULLSEL)
));
ap_MP2_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_7_PULLEN),
  .pullsel(`MP2_7_PULLSEL),
  .pad_pd(`MP2_7)
));
ap_MP2_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_7),
  .pullen(`MP2_7_PULLEN),
  .pullsel(`MP2_7_PULLSEL)
));
ap_MP2_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_8_OUTFUNC_SEL),
  .gpioouten(`MP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0TX_OE),
  .od(`MP2_8_PINCTRL_0_OD),
  .func_out(`LPD_LIN0TX_OUT),
  .pad(`MP2_8)
));
ap_MP2_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_8_OUTFUNC_SEL),
  .gpioouten(`MP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0TX_OE),
  .od(`MP2_8_PINCTRL_0_OD),
  .func_out(`LPD_LIN0TX_OUT),
  .pad(`MP2_8),
  .pad_gz(`MP2_8_pad_y)
));
ap_MP2_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_8_OUTFUNC_SEL),
  .gpioouten(`MP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`MP2_8_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`MP2_8)
));
ap_MP2_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_8_OUTFUNC_SEL),
  .gpioouten(`MP2_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4TX_OE),
  .od(`MP2_8_PINCTRL_0_OD),
  .func_out(`CAN4TX_OUT),
  .pad(`MP2_8),
  .pad_gz(`MP2_8_pad_y)
));
ap_MP2_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_8_PULLEN),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_8)
));
ap_MP2_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_8),
  .pullen(`MP2_8_PULLEN),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE)
));
ap_MP2_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_8_PINCTRL_0_IE),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_8),
  .pad(`MP2_8),
  .default_value(`default_value)));
ap_MP2_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_8_PULLEN),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_8)
));
ap_MP2_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_8),
  .pullen(`MP2_8_PULLEN),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE)
));
ap_MP2_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_8_PINCTRL_0_IE),
  .outen(`MP2_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_8),
  .pad(`MP2_8),
  .default_value(`default_value)));
ap_MP2_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_8_PULLEN),
  .pullsel(`MP2_8_PULLSEL),
  .pad_pullup(`MP2_8)
));
ap_MP2_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_8),
  .pullen(`MP2_8_PULLEN),
  .pullsel(`MP2_8_PULLSEL)
));
ap_MP2_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_8_PULLEN),
  .pullsel(`MP2_8_PULLSEL),
  .pad_pd(`MP2_8)
));
ap_MP2_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_8),
  .pullen(`MP2_8_PULLEN),
  .pullsel(`MP2_8_PULLSEL)
));
ap_MP2_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0RX_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`LPD_LIN0RX_OUT),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0RX_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`LPD_LIN0RX_OUT),
  .pad(`MP2_9),
  .pad_gz(`MP2_9_pad_y)
));
ap_MP2_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN4RX_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`CAN4RX_OUT),
  .pad(`MP2_9),
  .pad_gz(`MP2_9_pad_y)
));
ap_MP2_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_9),
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE)
));
ap_MP2_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_9_PINCTRL_0_IE),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_9),
  .pad(`MP2_9),
  .default_value(`default_value)));
ap_MP2_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_9),
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE)
));
ap_MP2_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_9_PINCTRL_0_IE),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_9),
  .pad(`MP2_9),
  .default_value(`default_value)));
ap_MP2_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_9_OUTFUNC_SEL),
  .gpioouten(`MP2_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS0_OE),
  .od(`MP2_9_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS0_OUT),
  .pad(`MP2_9),
  .pad_gz(`MP2_9_pad_y)
));
ap_MP2_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_9)
));
ap_MP2_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_9),
  .pullen(`MP2_9_PULLEN),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE)
));
ap_MP2_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_9_PINCTRL_0_IE),
  .outen(`MP2_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_9),
  .pad(`MP2_9),
  .default_value(`default_value)));
ap_MP2_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_9_PULLEN),
  .pullsel(`MP2_9_PULLSEL),
  .pad_pullup(`MP2_9)
));
ap_MP2_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_9),
  .pullen(`MP2_9_PULLEN),
  .pullsel(`MP2_9_PULLSEL)
));
ap_MP2_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_9_PULLEN),
  .pullsel(`MP2_9_PULLSEL),
  .pad_pd(`MP2_9)
));
ap_MP2_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_9),
  .pullen(`MP2_9_PULLEN),
  .pullsel(`MP2_9_PULLSEL)
));
ap_MP2_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP2_10),
  .pad_gz(`MP2_10_pad_y)
));
ap_MP2_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE)
));
ap_MP2_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_10_PINCTRL_0_IE),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_10),
  .pad(`MP2_10),
  .default_value(`default_value)));
ap_MP2_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5TX_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`CAN5TX_OUT),
  .pad(`MP2_10),
  .pad_gz(`MP2_10_pad_y)
));
ap_MP2_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE)
));
ap_MP2_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_10_PINCTRL_0_IE),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_10),
  .pad(`MP2_10),
  .default_value(`default_value)));
ap_MP2_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE)
));
ap_MP2_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_10_PINCTRL_0_IE),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_10),
  .pad(`MP2_10),
  .default_value(`default_value)));
ap_MP2_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_10_OUTFUNC_SEL),
  .gpioouten(`MP2_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS1_OE),
  .od(`MP2_10_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS1_OUT),
  .pad(`MP2_10),
  .pad_gz(`MP2_10_pad_y)
));
ap_MP2_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_10)
));
ap_MP2_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE)
));
ap_MP2_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_10_PINCTRL_0_IE),
  .outen(`MP2_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_10),
  .pad(`MP2_10),
  .default_value(`default_value)));
ap_MP2_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_10_PULLEN),
  .pullsel(`MP2_10_PULLSEL),
  .pad_pullup(`MP2_10)
));
ap_MP2_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .pullsel(`MP2_10_PULLSEL)
));
ap_MP2_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_10_PULLEN),
  .pullsel(`MP2_10_PULLSEL),
  .pad_pd(`MP2_10)
));
ap_MP2_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_10),
  .pullen(`MP2_10_PULLEN),
  .pullsel(`MP2_10_PULLSEL)
));
ap_MP2_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP2_11),
  .pad_gz(`MP2_11_pad_y)
));
ap_MP2_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE)
));
ap_MP2_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_11_PINCTRL_0_IE),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_11),
  .pad(`MP2_11),
  .default_value(`default_value)));
ap_MP2_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN5RX_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`CAN5RX_OUT),
  .pad(`MP2_11),
  .pad_gz(`MP2_11_pad_y)
));
ap_MP2_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE)
));
ap_MP2_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_11_PINCTRL_0_IE),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_11),
  .pad(`MP2_11),
  .default_value(`default_value)));
ap_MP2_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE)
));
ap_MP2_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_11_PINCTRL_0_IE),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_11),
  .pad(`MP2_11),
  .default_value(`default_value)));
ap_MP2_11_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_11_OUTFUNC_SEL),
  .gpioouten(`MP2_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS2_OE),
  .od(`MP2_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS2_OUT),
  .pad(`MP2_11),
  .pad_gz(`MP2_11_pad_y)
));
ap_MP2_11_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_11)
));
ap_MP2_11_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE)
));
ap_MP2_11_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_11_PINCTRL_0_IE),
  .outen(`MP2_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_11),
  .pad(`MP2_11),
  .default_value(`default_value)));
ap_MP2_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_11_PULLEN),
  .pullsel(`MP2_11_PULLSEL),
  .pad_pullup(`MP2_11)
));
ap_MP2_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .pullsel(`MP2_11_PULLSEL)
));
ap_MP2_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_11_PULLEN),
  .pullsel(`MP2_11_PULLSEL),
  .pad_pd(`MP2_11)
));
ap_MP2_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_11),
  .pullen(`MP2_11_PULLEN),
  .pullsel(`MP2_11_PULLSEL)
));
ap_MP2_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP2_12),
  .pad_gz(`MP2_12_pad_y)
));
ap_MP2_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE)
));
ap_MP2_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_12_PINCTRL_0_IE),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_12),
  .pad(`MP2_12),
  .default_value(`default_value)));
ap_MP2_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`MP2_12),
  .pad_gz(`MP2_12_pad_y)
));
ap_MP2_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE)
));
ap_MP2_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_12_PINCTRL_0_IE),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_12),
  .pad(`MP2_12),
  .default_value(`default_value)));
ap_MP2_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE)
));
ap_MP2_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_12_PINCTRL_0_IE),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_12),
  .pad(`MP2_12),
  .default_value(`default_value)));
ap_MP2_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_12_OUTFUNC_SEL),
  .gpioouten(`MP2_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS3_OE),
  .od(`MP2_12_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS3_OUT),
  .pad(`MP2_12),
  .pad_gz(`MP2_12_pad_y)
));
ap_MP2_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_12)
));
ap_MP2_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE)
));
ap_MP2_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_12_PINCTRL_0_IE),
  .outen(`MP2_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_12),
  .pad(`MP2_12),
  .default_value(`default_value)));
ap_MP2_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_12_PULLEN),
  .pullsel(`MP2_12_PULLSEL),
  .pad_pullup(`MP2_12)
));
ap_MP2_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .pullsel(`MP2_12_PULLSEL)
));
ap_MP2_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_12_PULLEN),
  .pullsel(`MP2_12_PULLSEL),
  .pad_pd(`MP2_12)
));
ap_MP2_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_12),
  .pullen(`MP2_12_PULLEN),
  .pullsel(`MP2_12_PULLSEL)
));
ap_MP2_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP2_13),
  .pad_gz(`MP2_13_pad_y)
));
ap_MP2_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE)
));
ap_MP2_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP2_13_PINCTRL_0_IE),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_13),
  .pad(`MP2_13),
  .default_value(`default_value)));
ap_MP2_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`MP2_13),
  .pad_gz(`MP2_13_pad_y)
));
ap_MP2_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE)
));
ap_MP2_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_13_PINCTRL_0_IE),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_13),
  .pad(`MP2_13),
  .default_value(`default_value)));
ap_MP2_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE)
));
ap_MP2_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_13_PINCTRL_0_IE),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_13),
  .pad(`MP2_13),
  .default_value(`default_value)));
ap_MP2_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_13_OUTFUNC_SEL),
  .gpioouten(`MP2_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP2_13_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP2_13),
  .pad_gz(`MP2_13_pad_y)
));
ap_MP2_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_13)
));
ap_MP2_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE)
));
ap_MP2_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_13_PINCTRL_0_IE),
  .outen(`MP2_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_13),
  .pad(`MP2_13),
  .default_value(`default_value)));
ap_MP2_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_13_PULLEN),
  .pullsel(`MP2_13_PULLSEL),
  .pad_pullup(`MP2_13)
));
ap_MP2_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .pullsel(`MP2_13_PULLSEL)
));
ap_MP2_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_13_PULLEN),
  .pullsel(`MP2_13_PULLSEL),
  .pad_pd(`MP2_13)
));
ap_MP2_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_13),
  .pullen(`MP2_13_PULLEN),
  .pullsel(`MP2_13_PULLSEL)
));
ap_MP2_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0TX_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`LPD_LIN0TX_OUT),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0TX_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`LPD_LIN0TX_OUT),
  .pad(`MP2_14),
  .pad_gz(`MP2_14_pad_y)
));
ap_MP2_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`MP2_14),
  .pad_gz(`MP2_14_pad_y)
));
ap_MP2_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_14),
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE)
));
ap_MP2_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_14_PINCTRL_0_IE),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_14),
  .pad(`MP2_14),
  .default_value(`default_value)));
ap_MP2_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_14),
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE)
));
ap_MP2_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_14_PINCTRL_0_IE),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_14),
  .pad(`MP2_14),
  .default_value(`default_value)));
ap_MP2_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_14_OUTFUNC_SEL),
  .gpioouten(`MP2_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP2_14_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP2_14),
  .pad_gz(`MP2_14_pad_y)
));
ap_MP2_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_14)
));
ap_MP2_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_14),
  .pullen(`MP2_14_PULLEN),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE)
));
ap_MP2_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_14_PINCTRL_0_IE),
  .outen(`MP2_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_14),
  .pad(`MP2_14),
  .default_value(`default_value)));
ap_MP2_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_14_PULLEN),
  .pullsel(`MP2_14_PULLSEL),
  .pad_pullup(`MP2_14)
));
ap_MP2_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_14),
  .pullen(`MP2_14_PULLEN),
  .pullsel(`MP2_14_PULLSEL)
));
ap_MP2_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_14_PULLEN),
  .pullsel(`MP2_14_PULLSEL),
  .pad_pd(`MP2_14)
));
ap_MP2_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_14),
  .pullen(`MP2_14_PULLEN),
  .pullsel(`MP2_14_PULLSEL)
));
ap_MP2_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0RX_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`LPD_LIN0RX_OUT),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`LPD_LIN0RX_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`LPD_LIN0RX_OUT),
  .pad(`MP2_15),
  .pad_gz(`MP2_15_pad_y)
));
ap_MP2_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`MP2_15),
  .pad_gz(`MP2_15_pad_y)
));
ap_MP2_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_15),
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE)
));
ap_MP2_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP2_15_PINCTRL_0_IE),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_15),
  .pad(`MP2_15),
  .default_value(`default_value)));
ap_MP2_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_15),
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE)
));
ap_MP2_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP2_15_PINCTRL_0_IE),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_15),
  .pad(`MP2_15),
  .default_value(`default_value)));
ap_MP2_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP2_15_OUTFUNC_SEL),
  .gpioouten(`MP2_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP2_15_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP2_15),
  .pad_gz(`MP2_15_pad_y)
));
ap_MP2_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP2_15)
));
ap_MP2_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP2_15),
  .pullen(`MP2_15_PULLEN),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE)
));
ap_MP2_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP2_15_PINCTRL_0_IE),
  .outen(`MP2_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP2_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP2_15),
  .pad(`MP2_15),
  .default_value(`default_value)));
ap_MP2_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP2_15_PULLEN),
  .pullsel(`MP2_15_PULLSEL),
  .pad_pullup(`MP2_15)
));
ap_MP2_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP2_15),
  .pullen(`MP2_15_PULLEN),
  .pullsel(`MP2_15_PULLSEL)
));
ap_MP2_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP2_15_PULLEN),
  .pullsel(`MP2_15_PULLSEL),
  .pad_pd(`MP2_15)
));
ap_MP2_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP2_15),
  .pullen(`MP2_15_PULLEN),
  .pullsel(`MP2_15_PULLSEL)
));
ap_MP0_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE)
));
ap_MP0_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_0_PINCTRL_0_IE),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_0),
  .pad(`MP0_0),
  .default_value(`default_value)));
ap_MP0_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`MP0_0),
  .pad_gz(`MP0_0_pad_y)
));
ap_MP0_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE)
));
ap_MP0_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_0_PINCTRL_0_IE),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_0),
  .pad(`MP0_0),
  .default_value(`default_value)));
ap_MP0_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP0_0),
  .pad_gz(`MP0_0_pad_y)
));
ap_MP0_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE)
));
ap_MP0_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_0_PINCTRL_0_IE),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_0),
  .pad(`MP0_0),
  .default_value(`default_value)));
ap_MP0_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_0_OUTFUNC_SEL),
  .gpioouten(`MP0_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP0_0_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP0_0),
  .pad_gz(`MP0_0_pad_y)
));
ap_MP0_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_0)
));
ap_MP0_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE)
));
ap_MP0_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_0_PINCTRL_0_IE),
  .outen(`MP0_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_0),
  .pad(`MP0_0),
  .default_value(`default_value)));
ap_MP0_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_0_PULLEN),
  .pullsel(`MP0_0_PULLSEL),
  .pad_pullup(`MP0_0)
));
ap_MP0_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .pullsel(`MP0_0_PULLSEL)
));
ap_MP0_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_0_PULLEN),
  .pullsel(`MP0_0_PULLSEL),
  .pad_pd(`MP0_0)
));
ap_MP0_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_0),
  .pullen(`MP0_0_PULLEN),
  .pullsel(`MP0_0_PULLSEL)
));
ap_MP0_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE)
));
ap_MP0_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_1_PINCTRL_0_IE),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_1),
  .pad(`MP0_1),
  .default_value(`default_value)));
ap_MP0_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`MP0_1),
  .pad_gz(`MP0_1_pad_y)
));
ap_MP0_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE)
));
ap_MP0_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_1_PINCTRL_0_IE),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_1),
  .pad(`MP0_1),
  .default_value(`default_value)));
ap_MP0_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP0_1),
  .pad_gz(`MP0_1_pad_y)
));
ap_MP0_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE)
));
ap_MP0_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_1_PINCTRL_0_IE),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_1),
  .pad(`MP0_1),
  .default_value(`default_value)));
ap_MP0_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_1_OUTFUNC_SEL),
  .gpioouten(`MP0_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP0_1_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP0_1),
  .pad_gz(`MP0_1_pad_y)
));
ap_MP0_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_1)
));
ap_MP0_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE)
));
ap_MP0_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_1_PINCTRL_0_IE),
  .outen(`MP0_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_1),
  .pad(`MP0_1),
  .default_value(`default_value)));
ap_MP0_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_1_PULLEN),
  .pullsel(`MP0_1_PULLSEL),
  .pad_pullup(`MP0_1)
));
ap_MP0_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .pullsel(`MP0_1_PULLSEL)
));
ap_MP0_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_1_PULLEN),
  .pullsel(`MP0_1_PULLSEL),
  .pad_pd(`MP0_1)
));
ap_MP0_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_1),
  .pullen(`MP0_1_PULLEN),
  .pullsel(`MP0_1_PULLSEL)
));
ap_MP0_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE)
));
ap_MP0_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_2_PINCTRL_0_IE),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_2),
  .pad(`MP0_2),
  .default_value(`default_value)));
ap_MP0_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`MP0_2),
  .pad_gz(`MP0_2_pad_y)
));
ap_MP0_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE)
));
ap_MP0_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_2_PINCTRL_0_IE),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_2),
  .pad(`MP0_2),
  .default_value(`default_value)));
ap_MP0_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP0_2),
  .pad_gz(`MP0_2_pad_y)
));
ap_MP0_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE)
));
ap_MP0_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_2_PINCTRL_0_IE),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_2),
  .pad(`MP0_2),
  .default_value(`default_value)));
ap_MP0_2_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_2_OUTFUNC_SEL),
  .gpioouten(`MP0_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP0_2_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP0_2),
  .pad_gz(`MP0_2_pad_y)
));
ap_MP0_2_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_2)
));
ap_MP0_2_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE)
));
ap_MP0_2_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_2_PINCTRL_0_IE),
  .outen(`MP0_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_2),
  .pad(`MP0_2),
  .default_value(`default_value)));
ap_MP0_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_2_PULLEN),
  .pullsel(`MP0_2_PULLSEL),
  .pad_pullup(`MP0_2)
));
ap_MP0_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .pullsel(`MP0_2_PULLSEL)
));
ap_MP0_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_2_PULLEN),
  .pullsel(`MP0_2_PULLSEL),
  .pad_pd(`MP0_2)
));
ap_MP0_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_2),
  .pullen(`MP0_2_PULLEN),
  .pullsel(`MP0_2_PULLSEL)
));
ap_MP0_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE)
));
ap_MP0_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_3_PINCTRL_0_IE),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_3),
  .pad(`MP0_3),
  .default_value(`default_value)));
ap_MP0_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`MP0_3),
  .pad_gz(`MP0_3_pad_y)
));
ap_MP0_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE)
));
ap_MP0_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_3_PINCTRL_0_IE),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_3),
  .pad(`MP0_3),
  .default_value(`default_value)));
ap_MP0_3_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP0_3),
  .pad_gz(`MP0_3_pad_y)
));
ap_MP0_3_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE)
));
ap_MP0_3_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_3_PINCTRL_0_IE),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_3),
  .pad(`MP0_3),
  .default_value(`default_value)));
ap_MP0_3_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_3_OUTFUNC_SEL),
  .gpioouten(`MP0_3_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP0_3_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP0_3),
  .pad_gz(`MP0_3_pad_y)
));
ap_MP0_3_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_3)
));
ap_MP0_3_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE)
));
ap_MP0_3_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_3_PINCTRL_0_IE),
  .outen(`MP0_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_3),
  .pad(`MP0_3),
  .default_value(`default_value)));
ap_MP0_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_3_PULLEN),
  .pullsel(`MP0_3_PULLSEL),
  .pad_pullup(`MP0_3)
));
ap_MP0_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .pullsel(`MP0_3_PULLSEL)
));
ap_MP0_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_3_PULLEN),
  .pullsel(`MP0_3_PULLSEL),
  .pad_pd(`MP0_3)
));
ap_MP0_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_3),
  .pullen(`MP0_3_PULLEN),
  .pullsel(`MP0_3_PULLSEL)
));
ap_MP0_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE)
));
ap_MP0_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_4_PINCTRL_0_IE),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_4),
  .pad(`MP0_4),
  .default_value(`default_value)));
ap_MP0_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`MP0_4),
  .pad_gz(`MP0_4_pad_y)
));
ap_MP0_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE)
));
ap_MP0_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_4_PINCTRL_0_IE),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_4),
  .pad(`MP0_4),
  .default_value(`default_value)));
ap_MP0_4_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP0_4),
  .pad_gz(`MP0_4_pad_y)
));
ap_MP0_4_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE)
));
ap_MP0_4_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_4_PINCTRL_0_IE),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_4),
  .pad(`MP0_4),
  .default_value(`default_value)));
ap_MP0_4_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_4_OUTFUNC_SEL),
  .gpioouten(`MP0_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP0_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP0_4),
  .pad_gz(`MP0_4_pad_y)
));
ap_MP0_4_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_4)
));
ap_MP0_4_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE)
));
ap_MP0_4_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_4_PINCTRL_0_IE),
  .outen(`MP0_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_4),
  .pad(`MP0_4),
  .default_value(`default_value)));
ap_MP0_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_4_PULLEN),
  .pullsel(`MP0_4_PULLSEL),
  .pad_pullup(`MP0_4)
));
ap_MP0_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .pullsel(`MP0_4_PULLSEL)
));
ap_MP0_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_4_PULLEN),
  .pullsel(`MP0_4_PULLSEL),
  .pad_pd(`MP0_4)
));
ap_MP0_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_4),
  .pullen(`MP0_4_PULLEN),
  .pullsel(`MP0_4_PULLSEL)
));
ap_MP0_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_5_PULLEN),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_5)
));
ap_MP0_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_5),
  .pullen(`MP0_5_PULLEN),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE)
));
ap_MP0_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_5_PINCTRL_0_IE),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_5),
  .pad(`MP0_5),
  .default_value(`default_value)));
ap_MP0_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_5_OUTFUNC_SEL),
  .gpioouten(`MP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`MP0_5_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`MP0_5)
));
ap_MP0_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_5_OUTFUNC_SEL),
  .gpioouten(`MP0_5_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`MP0_5_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`MP0_5),
  .pad_gz(`MP0_5_pad_y)
));
ap_MP0_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_5_PULLEN),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_5)
));
ap_MP0_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_5),
  .pullen(`MP0_5_PULLEN),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE)
));
ap_MP0_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_5_PINCTRL_0_IE),
  .outen(`MP0_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_5),
  .pad(`MP0_5),
  .default_value(`default_value)));
ap_MP0_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_5_PULLEN),
  .pullsel(`MP0_5_PULLSEL),
  .pad_pullup(`MP0_5)
));
ap_MP0_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_5),
  .pullen(`MP0_5_PULLEN),
  .pullsel(`MP0_5_PULLSEL)
));
ap_MP0_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_5_PULLEN),
  .pullsel(`MP0_5_PULLSEL),
  .pad_pd(`MP0_5)
));
ap_MP0_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_5),
  .pullen(`MP0_5_PULLEN),
  .pullsel(`MP0_5_PULLSEL)
));
ap_MP0_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE)
));
ap_MP0_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_6_PINCTRL_0_IE),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_6),
  .pad(`MP0_6),
  .default_value(`default_value)));
ap_MP0_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP0_6),
  .pad_gz(`MP0_6_pad_y)
));
ap_MP0_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE)
));
ap_MP0_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_6_PINCTRL_0_IE),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_6),
  .pad(`MP0_6),
  .default_value(`default_value)));
ap_MP0_6_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP0_6),
  .pad_gz(`MP0_6_pad_y)
));
ap_MP0_6_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE)
));
ap_MP0_6_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_6_PINCTRL_0_IE),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_6),
  .pad(`MP0_6),
  .default_value(`default_value)));
ap_MP0_6_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_6_OUTFUNC_SEL),
  .gpioouten(`MP0_6_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS4_OE),
  .od(`MP0_6_PINCTRL_0_OD),
  .func_out(`SPI8CS4_OUT),
  .pad(`MP0_6),
  .pad_gz(`MP0_6_pad_y)
));
ap_MP0_6_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_6)
));
ap_MP0_6_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE)
));
ap_MP0_6_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_6_PINCTRL_0_IE),
  .outen(`MP0_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_6),
  .pad(`MP0_6),
  .default_value(`default_value)));
ap_MP0_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_6_PULLEN),
  .pullsel(`MP0_6_PULLSEL),
  .pad_pullup(`MP0_6)
));
ap_MP0_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .pullsel(`MP0_6_PULLSEL)
));
ap_MP0_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_6_PULLEN),
  .pullsel(`MP0_6_PULLSEL),
  .pad_pd(`MP0_6)
));
ap_MP0_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_6),
  .pullen(`MP0_6_PULLEN),
  .pullsel(`MP0_6_PULLSEL)
));
ap_MP0_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE)
));
ap_MP0_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_7_PINCTRL_0_IE),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_7),
  .pad(`MP0_7),
  .default_value(`default_value)));
ap_MP0_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP0_7),
  .pad_gz(`MP0_7_pad_y)
));
ap_MP0_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE)
));
ap_MP0_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_7_PINCTRL_0_IE),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_7),
  .pad(`MP0_7),
  .default_value(`default_value)));
ap_MP0_7_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP0_7),
  .pad_gz(`MP0_7_pad_y)
));
ap_MP0_7_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE)
));
ap_MP0_7_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_7_PINCTRL_0_IE),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_7),
  .pad(`MP0_7),
  .default_value(`default_value)));
ap_MP0_7_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_7_OUTFUNC_SEL),
  .gpioouten(`MP0_7_GPIO_OUTPUT_ENABLE),
  .oe(`SPI8CS5_OE),
  .od(`MP0_7_PINCTRL_0_OD),
  .func_out(`SPI8CS5_OUT),
  .pad(`MP0_7),
  .pad_gz(`MP0_7_pad_y)
));
ap_MP0_7_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_7)
));
ap_MP0_7_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE)
));
ap_MP0_7_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_7_PINCTRL_0_IE),
  .outen(`MP0_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_7),
  .pad(`MP0_7),
  .default_value(`default_value)));
ap_MP0_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_7_PULLEN),
  .pullsel(`MP0_7_PULLSEL),
  .pad_pullup(`MP0_7)
));
ap_MP0_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .pullsel(`MP0_7_PULLSEL)
));
ap_MP0_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_7_PULLEN),
  .pullsel(`MP0_7_PULLSEL),
  .pad_pd(`MP0_7)
));
ap_MP0_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_7),
  .pullen(`MP0_7_PULLEN),
  .pullsel(`MP0_7_PULLSEL)
));
ap_MP0_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6TX_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`CAN6TX_OUT),
  .pad(`MP0_8),
  .pad_gz(`MP0_8_pad_y)
));
ap_MP0_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE)
));
ap_MP0_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_8_PINCTRL_0_IE),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_8),
  .pad(`MP0_8),
  .default_value(`default_value)));
ap_MP0_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0TX_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`LIN0TX_OUT),
  .pad(`MP0_8),
  .pad_gz(`MP0_8_pad_y)
));
ap_MP0_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE)
));
ap_MP0_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_8_PINCTRL_0_IE),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_8),
  .pad(`MP0_8),
  .default_value(`default_value)));
ap_MP0_8_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE)
));
ap_MP0_8_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_8_PINCTRL_0_IE),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_8),
  .pad(`MP0_8),
  .default_value(`default_value)));
ap_MP0_8_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP0_8),
  .pad_gz(`MP0_8_pad_y)
));
ap_MP0_8_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE)
));
ap_MP0_8_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_8_PINCTRL_0_IE),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_8),
  .pad(`MP0_8),
  .default_value(`default_value)));
ap_MP0_8_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_8_OUTFUNC_SEL),
  .gpioouten(`MP0_8_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS4_OE),
  .od(`MP0_8_PINCTRL_0_OD),
  .func_out(`SPI9CS4_OUT),
  .pad(`MP0_8),
  .pad_gz(`MP0_8_pad_y)
));
ap_MP0_8_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_8)
));
ap_MP0_8_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE)
));
ap_MP0_8_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP0_8_PINCTRL_0_IE),
  .outen(`MP0_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_8),
  .pad(`MP0_8),
  .default_value(`default_value)));
ap_MP0_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_8_PULLEN),
  .pullsel(`MP0_8_PULLSEL),
  .pad_pullup(`MP0_8)
));
ap_MP0_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .pullsel(`MP0_8_PULLSEL)
));
ap_MP0_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_8_PULLEN),
  .pullsel(`MP0_8_PULLSEL),
  .pad_pd(`MP0_8)
));
ap_MP0_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_8),
  .pullen(`MP0_8_PULLEN),
  .pullsel(`MP0_8_PULLSEL)
));
ap_MP0_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`CAN6RX_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`CAN6RX_OUT),
  .pad(`MP0_9),
  .pad_gz(`MP0_9_pad_y)
));
ap_MP0_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE)
));
ap_MP0_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_9_PINCTRL_0_IE),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_9),
  .pad(`MP0_9),
  .default_value(`default_value)));
ap_MP0_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`LIN0RX_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`LIN0RX_OUT),
  .pad(`MP0_9),
  .pad_gz(`MP0_9_pad_y)
));
ap_MP0_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE)
));
ap_MP0_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_9_PINCTRL_0_IE),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_9),
  .pad(`MP0_9),
  .default_value(`default_value)));
ap_MP0_9_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE)
));
ap_MP0_9_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_9_PINCTRL_0_IE),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_9),
  .pad(`MP0_9),
  .default_value(`default_value)));
ap_MP0_9_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_9_OUTFUNC_SEL),
  .gpioouten(`MP0_9_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP0_9_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP0_9),
  .pad_gz(`MP0_9_pad_y)
));
ap_MP0_9_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_9)
));
ap_MP0_9_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE)
));
ap_MP0_9_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_9_PINCTRL_0_IE),
  .outen(`MP0_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_9),
  .pad(`MP0_9),
  .default_value(`default_value)));
ap_MP0_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_9_PULLEN),
  .pullsel(`MP0_9_PULLSEL),
  .pad_pullup(`MP0_9)
));
ap_MP0_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .pullsel(`MP0_9_PULLSEL)
));
ap_MP0_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_9_PULLEN),
  .pullsel(`MP0_9_PULLSEL),
  .pad_pd(`MP0_9)
));
ap_MP0_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_9),
  .pullen(`MP0_9_PULLEN),
  .pullsel(`MP0_9_PULLSEL)
));
ap_MP0_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7TX_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`CAN7TX_OUT),
  .pad(`MP0_10),
  .pad_gz(`MP0_10_pad_y)
));
ap_MP0_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE)
));
ap_MP0_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_10_PINCTRL_0_IE),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_10),
  .pad(`MP0_10),
  .default_value(`default_value)));
ap_MP0_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`MP0_10),
  .pad_gz(`MP0_10_pad_y)
));
ap_MP0_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE)
));
ap_MP0_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_10_PINCTRL_0_IE),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_10),
  .pad(`MP0_10),
  .default_value(`default_value)));
ap_MP0_10_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE)
));
ap_MP0_10_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_10_PINCTRL_0_IE),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_10),
  .pad(`MP0_10),
  .default_value(`default_value)));
ap_MP0_10_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_10_OUTFUNC_SEL),
  .gpioouten(`MP0_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP0_10_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP0_10),
  .pad_gz(`MP0_10_pad_y)
));
ap_MP0_10_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_10)
));
ap_MP0_10_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE)
));
ap_MP0_10_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_10_PINCTRL_0_IE),
  .outen(`MP0_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_10),
  .pad(`MP0_10),
  .default_value(`default_value)));
ap_MP0_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_10_PULLEN),
  .pullsel(`MP0_10_PULLSEL),
  .pad_pullup(`MP0_10)
));
ap_MP0_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .pullsel(`MP0_10_PULLSEL)
));
ap_MP0_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_10_PULLEN),
  .pullsel(`MP0_10_PULLSEL),
  .pad_pd(`MP0_10)
));
ap_MP0_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_10),
  .pullen(`MP0_10_PULLEN),
  .pullsel(`MP0_10_PULLSEL)
));
ap_MP0_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_11_OUTFUNC_SEL),
  .gpioouten(`MP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`MP0_11_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`MP0_11)
));
ap_MP0_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_11_OUTFUNC_SEL),
  .gpioouten(`MP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`CAN7RX_OE),
  .od(`MP0_11_PINCTRL_0_OD),
  .func_out(`CAN7RX_OUT),
  .pad(`MP0_11),
  .pad_gz(`MP0_11_pad_y)
));
ap_MP0_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_11)
));
ap_MP0_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_11),
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE)
));
ap_MP0_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_11_PINCTRL_0_IE),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_11),
  .pad(`MP0_11),
  .default_value(`default_value)));
ap_MP0_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_11_OUTFUNC_SEL),
  .gpioouten(`MP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`MP0_11_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`MP0_11)
));
ap_MP0_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_11_OUTFUNC_SEL),
  .gpioouten(`MP0_11_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`MP0_11_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`MP0_11),
  .pad_gz(`MP0_11_pad_y)
));
ap_MP0_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_11)
));
ap_MP0_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_11),
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE)
));
ap_MP0_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_11_PINCTRL_0_IE),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_11),
  .pad(`MP0_11),
  .default_value(`default_value)));
ap_MP0_11_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_11)
));
ap_MP0_11_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_11),
  .pullen(`MP0_11_PULLEN),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE)
));
ap_MP0_11_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_11_PINCTRL_0_IE),
  .outen(`MP0_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_11),
  .pad(`MP0_11),
  .default_value(`default_value)));
ap_MP0_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_11_PULLEN),
  .pullsel(`MP0_11_PULLSEL),
  .pad_pullup(`MP0_11)
));
ap_MP0_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_11),
  .pullen(`MP0_11_PULLEN),
  .pullsel(`MP0_11_PULLSEL)
));
ap_MP0_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_11_PULLEN),
  .pullsel(`MP0_11_PULLSEL),
  .pad_pd(`MP0_11)
));
ap_MP0_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_11),
  .pullen(`MP0_11_PULLEN),
  .pullsel(`MP0_11_PULLSEL)
));
ap_MP0_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8TX_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`CAN8TX_OUT),
  .pad(`MP0_12),
  .pad_gz(`MP0_12_pad_y)
));
ap_MP0_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE)
));
ap_MP0_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_12_PINCTRL_0_IE),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_12),
  .pad(`MP0_12),
  .default_value(`default_value)));
ap_MP0_12_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2TX_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`LIN2TX_OUT),
  .pad(`MP0_12),
  .pad_gz(`MP0_12_pad_y)
));
ap_MP0_12_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE)
));
ap_MP0_12_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_12_PINCTRL_0_IE),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_12),
  .pad(`MP0_12),
  .default_value(`default_value)));
ap_MP0_12_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE)
));
ap_MP0_12_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_12_PINCTRL_0_IE),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_12),
  .pad(`MP0_12),
  .default_value(`default_value)));
ap_MP0_12_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_12_OUTFUNC_SEL),
  .gpioouten(`MP0_12_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`MP0_12_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`MP0_12),
  .pad_gz(`MP0_12_pad_y)
));
ap_MP0_12_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_12)
));
ap_MP0_12_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE)
));
ap_MP0_12_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_12_PINCTRL_0_IE),
  .outen(`MP0_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_12),
  .pad(`MP0_12),
  .default_value(`default_value)));
ap_MP0_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_12_PULLEN),
  .pullsel(`MP0_12_PULLSEL),
  .pad_pullup(`MP0_12)
));
ap_MP0_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .pullsel(`MP0_12_PULLSEL)
));
ap_MP0_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_12_PULLEN),
  .pullsel(`MP0_12_PULLSEL),
  .pad_pd(`MP0_12)
));
ap_MP0_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_12),
  .pullen(`MP0_12_PULLEN),
  .pullsel(`MP0_12_PULLSEL)
));
ap_MP0_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`CAN8RX_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`CAN8RX_OUT),
  .pad(`MP0_13),
  .pad_gz(`MP0_13_pad_y)
));
ap_MP0_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE)
));
ap_MP0_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_13_PINCTRL_0_IE),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_13),
  .pad(`MP0_13),
  .default_value(`default_value)));
ap_MP0_13_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`LIN2RX_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`LIN2RX_OUT),
  .pad(`MP0_13),
  .pad_gz(`MP0_13_pad_y)
));
ap_MP0_13_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE)
));
ap_MP0_13_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_13_PINCTRL_0_IE),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_13),
  .pad(`MP0_13),
  .default_value(`default_value)));
ap_MP0_13_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE)
));
ap_MP0_13_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_13_PINCTRL_0_IE),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_13),
  .pad(`MP0_13),
  .default_value(`default_value)));
ap_MP0_13_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_13_OUTFUNC_SEL),
  .gpioouten(`MP0_13_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`MP0_13_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`MP0_13),
  .pad_gz(`MP0_13_pad_y)
));
ap_MP0_13_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_13)
));
ap_MP0_13_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE)
));
ap_MP0_13_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_13_PINCTRL_0_IE),
  .outen(`MP0_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_13),
  .pad(`MP0_13),
  .default_value(`default_value)));
ap_MP0_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_13_PULLEN),
  .pullsel(`MP0_13_PULLSEL),
  .pad_pullup(`MP0_13)
));
ap_MP0_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .pullsel(`MP0_13_PULLSEL)
));
ap_MP0_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_13_PULLEN),
  .pullsel(`MP0_13_PULLSEL),
  .pad_pd(`MP0_13)
));
ap_MP0_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_13),
  .pullen(`MP0_13_PULLEN),
  .pullsel(`MP0_13_PULLSEL)
));
ap_MP0_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9TX_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`CAN9TX_OUT),
  .pad(`MP0_14),
  .pad_gz(`MP0_14_pad_y)
));
ap_MP0_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE)
));
ap_MP0_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_14_PINCTRL_0_IE),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_14),
  .pad(`MP0_14),
  .default_value(`default_value)));
ap_MP0_14_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS4_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`SPI3CS4_OUT),
  .pad(`MP0_14),
  .pad_gz(`MP0_14_pad_y)
));
ap_MP0_14_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE)
));
ap_MP0_14_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_14_PINCTRL_0_IE),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_14),
  .pad(`MP0_14),
  .default_value(`default_value)));
ap_MP0_14_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS4_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`SPI4CS4_OUT),
  .pad(`MP0_14),
  .pad_gz(`MP0_14_pad_y)
));
ap_MP0_14_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE)
));
ap_MP0_14_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_14_PINCTRL_0_IE),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_14),
  .pad(`MP0_14),
  .default_value(`default_value)));
ap_MP0_14_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_14_OUTFUNC_SEL),
  .gpioouten(`MP0_14_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1TX_OE),
  .od(`MP0_14_PINCTRL_0_OD),
  .func_out(`LIN1TX_OUT),
  .pad(`MP0_14),
  .pad_gz(`MP0_14_pad_y)
));
ap_MP0_14_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_14)
));
ap_MP0_14_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE)
));
ap_MP0_14_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_14_PINCTRL_0_IE),
  .outen(`MP0_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_14),
  .pad(`MP0_14),
  .default_value(`default_value)));
ap_MP0_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_14_PULLEN),
  .pullsel(`MP0_14_PULLSEL),
  .pad_pullup(`MP0_14)
));
ap_MP0_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .pullsel(`MP0_14_PULLSEL)
));
ap_MP0_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_14_PULLEN),
  .pullsel(`MP0_14_PULLSEL),
  .pad_pd(`MP0_14)
));
ap_MP0_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_14),
  .pullen(`MP0_14_PULLEN),
  .pullsel(`MP0_14_PULLSEL)
));
ap_MP0_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`CAN9RX_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`CAN9RX_OUT),
  .pad(`MP0_15),
  .pad_gz(`MP0_15_pad_y)
));
ap_MP0_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE)
));
ap_MP0_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_15_PINCTRL_0_IE),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_15),
  .pad(`MP0_15),
  .default_value(`default_value)));
ap_MP0_15_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI3CS5_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`SPI3CS5_OUT),
  .pad(`MP0_15),
  .pad_gz(`MP0_15_pad_y)
));
ap_MP0_15_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE)
));
ap_MP0_15_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_15_PINCTRL_0_IE),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_15),
  .pad(`MP0_15),
  .default_value(`default_value)));
ap_MP0_15_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`SPI4CS5_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`SPI4CS5_OUT),
  .pad(`MP0_15),
  .pad_gz(`MP0_15_pad_y)
));
ap_MP0_15_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE)
));
ap_MP0_15_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_15_PINCTRL_0_IE),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_15),
  .pad(`MP0_15),
  .default_value(`default_value)));
ap_MP0_15_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_15_OUTFUNC_SEL),
  .gpioouten(`MP0_15_GPIO_OUTPUT_ENABLE),
  .oe(`LIN1RX_OE),
  .od(`MP0_15_PINCTRL_0_OD),
  .func_out(`LIN1RX_OUT),
  .pad(`MP0_15),
  .pad_gz(`MP0_15_pad_y)
));
ap_MP0_15_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_15)
));
ap_MP0_15_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE)
));
ap_MP0_15_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_15_PINCTRL_0_IE),
  .outen(`MP0_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_15),
  .pad(`MP0_15),
  .default_value(`default_value)));
ap_MP0_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_15_PULLEN),
  .pullsel(`MP0_15_PULLSEL),
  .pad_pullup(`MP0_15)
));
ap_MP0_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .pullsel(`MP0_15_PULLSEL)
));
ap_MP0_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_15_PULLEN),
  .pullsel(`MP0_15_PULLSEL),
  .pad_pd(`MP0_15)
));
ap_MP0_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_15),
  .pullen(`MP0_15_PULLEN),
  .pullsel(`MP0_15_PULLSEL)
));
ap_MP0_16_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10TX_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`CAN10TX_OUT),
  .pad(`MP0_16),
  .pad_gz(`MP0_16_pad_y)
));
ap_MP0_16_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE)
));
ap_MP0_16_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_16_PINCTRL_0_IE),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_16),
  .pad(`MP0_16),
  .default_value(`default_value)));
ap_MP0_16_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`MP0_16),
  .pad_gz(`MP0_16_pad_y)
));
ap_MP0_16_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE)
));
ap_MP0_16_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_16_PINCTRL_0_IE),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_16),
  .pad(`MP0_16),
  .default_value(`default_value)));
ap_MP0_16_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS10_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS10_OUT),
  .pad(`MP0_16),
  .pad_gz(`MP0_16_pad_y)
));
ap_MP0_16_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE)
));
ap_MP0_16_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_16_PINCTRL_0_IE),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_16),
  .pad(`MP0_16),
  .default_value(`default_value)));
ap_MP0_16_FUNCSEL_5_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_5_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_16_OUTFUNC_SEL),
  .gpioouten(`MP0_16_GPIO_OUTPUT_ENABLE),
  .oe(`SPI9CS5_OE),
  .od(`MP0_16_PINCTRL_0_OD),
  .func_out(`SPI9CS5_OUT),
  .pad(`MP0_16),
  .pad_gz(`MP0_16_pad_y)
));
ap_MP0_16_FUNCSEL_5_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_16)
));
ap_MP0_16_FUNCSEL_5_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE)
));
ap_MP0_16_FUNCSEL_5_input_chk : assert property(iomux_input_path(
  .ie(`MP0_16_PINCTRL_0_IE),
  .outen(`MP0_16_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_16_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_16),
  .pad(`MP0_16),
  .default_value(`default_value)));
ap_MP0_16_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_16_PULLEN),
  .pullsel(`MP0_16_PULLSEL),
  .pad_pullup(`MP0_16)
));
ap_MP0_16_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .pullsel(`MP0_16_PULLSEL)
));
ap_MP0_16_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_16_PULLEN),
  .pullsel(`MP0_16_PULLSEL),
  .pad_pd(`MP0_16)
));
ap_MP0_16_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_16),
  .pullen(`MP0_16_PULLEN),
  .pullsel(`MP0_16_PULLSEL)
));
ap_MP0_17_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_17_OUTFUNC_SEL),
  .gpioouten(`MP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`MP0_17_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`MP0_17)
));
ap_MP0_17_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_17_OUTFUNC_SEL),
  .gpioouten(`MP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`CAN10RX_OE),
  .od(`MP0_17_PINCTRL_0_OD),
  .func_out(`CAN10RX_OUT),
  .pad(`MP0_17),
  .pad_gz(`MP0_17_pad_y)
));
ap_MP0_17_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_17_PULLEN),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_17)
));
ap_MP0_17_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_17),
  .pullen(`MP0_17_PULLEN),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE)
));
ap_MP0_17_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_17_PINCTRL_0_IE),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_17),
  .pad(`MP0_17),
  .default_value(`default_value)));
ap_MP0_17_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_17_OUTFUNC_SEL),
  .gpioouten(`MP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`MP0_17_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`MP0_17)
));
ap_MP0_17_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_17_OUTFUNC_SEL),
  .gpioouten(`MP0_17_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`MP0_17_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`MP0_17),
  .pad_gz(`MP0_17_pad_y)
));
ap_MP0_17_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_17_PULLEN),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_17)
));
ap_MP0_17_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_17),
  .pullen(`MP0_17_PULLEN),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE)
));
ap_MP0_17_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_17_PINCTRL_0_IE),
  .outen(`MP0_17_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_17_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_17),
  .pad(`MP0_17),
  .default_value(`default_value)));
ap_MP0_17_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_17_PULLEN),
  .pullsel(`MP0_17_PULLSEL),
  .pad_pullup(`MP0_17)
));
ap_MP0_17_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_17),
  .pullen(`MP0_17_PULLEN),
  .pullsel(`MP0_17_PULLSEL)
));
ap_MP0_17_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_17_PULLEN),
  .pullsel(`MP0_17_PULLSEL),
  .pad_pd(`MP0_17)
));
ap_MP0_17_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_17),
  .pullen(`MP0_17_PULLEN),
  .pullsel(`MP0_17_PULLSEL)
));
ap_MP0_18_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11TX_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`CAN11TX_OUT),
  .pad(`MP0_18),
  .pad_gz(`MP0_18_pad_y)
));
ap_MP0_18_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE)
));
ap_MP0_18_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_18_PINCTRL_0_IE),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_18),
  .pad(`MP0_18),
  .default_value(`default_value)));
ap_MP0_18_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`MP0_18),
  .pad_gz(`MP0_18_pad_y)
));
ap_MP0_18_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE)
));
ap_MP0_18_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_18_PINCTRL_0_IE),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_18),
  .pad(`MP0_18),
  .default_value(`default_value)));
ap_MP0_18_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS0_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS0_OUT),
  .pad(`MP0_18),
  .pad_gz(`MP0_18_pad_y)
));
ap_MP0_18_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE)
));
ap_MP0_18_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_18_PINCTRL_0_IE),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_18),
  .pad(`MP0_18),
  .default_value(`default_value)));
ap_MP0_18_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_18_OUTFUNC_SEL),
  .gpioouten(`MP0_18_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP0_18_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP0_18),
  .pad_gz(`MP0_18_pad_y)
));
ap_MP0_18_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_18)
));
ap_MP0_18_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE)
));
ap_MP0_18_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_18_PINCTRL_0_IE),
  .outen(`MP0_18_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_18_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_18),
  .pad(`MP0_18),
  .default_value(`default_value)));
ap_MP0_18_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_18_PULLEN),
  .pullsel(`MP0_18_PULLSEL),
  .pad_pullup(`MP0_18)
));
ap_MP0_18_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .pullsel(`MP0_18_PULLSEL)
));
ap_MP0_18_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_18_PULLEN),
  .pullsel(`MP0_18_PULLSEL),
  .pad_pd(`MP0_18)
));
ap_MP0_18_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_18),
  .pullen(`MP0_18_PULLEN),
  .pullsel(`MP0_18_PULLSEL)
));
ap_MP0_19_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`CAN11RX_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`CAN11RX_OUT),
  .pad(`MP0_19),
  .pad_gz(`MP0_19_pad_y)
));
ap_MP0_19_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE)
));
ap_MP0_19_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_19_PINCTRL_0_IE),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_19),
  .pad(`MP0_19),
  .default_value(`default_value)));
ap_MP0_19_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`MP0_19),
  .pad_gz(`MP0_19_pad_y)
));
ap_MP0_19_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE)
));
ap_MP0_19_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_19_PINCTRL_0_IE),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_19),
  .pad(`MP0_19),
  .default_value(`default_value)));
ap_MP0_19_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS1_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS1_OUT),
  .pad(`MP0_19),
  .pad_gz(`MP0_19_pad_y)
));
ap_MP0_19_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE)
));
ap_MP0_19_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_19_PINCTRL_0_IE),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_19),
  .pad(`MP0_19),
  .default_value(`default_value)));
ap_MP0_19_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_19_OUTFUNC_SEL),
  .gpioouten(`MP0_19_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP0_19_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP0_19),
  .pad_gz(`MP0_19_pad_y)
));
ap_MP0_19_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_19)
));
ap_MP0_19_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE)
));
ap_MP0_19_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_19_PINCTRL_0_IE),
  .outen(`MP0_19_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_19_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_19),
  .pad(`MP0_19),
  .default_value(`default_value)));
ap_MP0_19_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_19_PULLEN),
  .pullsel(`MP0_19_PULLSEL),
  .pad_pullup(`MP0_19)
));
ap_MP0_19_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .pullsel(`MP0_19_PULLSEL)
));
ap_MP0_19_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_19_PULLEN),
  .pullsel(`MP0_19_PULLSEL),
  .pad_pd(`MP0_19)
));
ap_MP0_19_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_19),
  .pullen(`MP0_19_PULLEN),
  .pullsel(`MP0_19_PULLSEL)
));
ap_MP0_20_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`MP0_20),
  .pad_gz(`MP0_20_pad_y)
));
ap_MP0_20_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE)
));
ap_MP0_20_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_20_PINCTRL_0_IE),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_20),
  .pad(`MP0_20),
  .default_value(`default_value)));
ap_MP0_20_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`MP0_20),
  .pad_gz(`MP0_20_pad_y)
));
ap_MP0_20_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE)
));
ap_MP0_20_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_20_PINCTRL_0_IE),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_20),
  .pad(`MP0_20),
  .default_value(`default_value)));
ap_MP0_20_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS2_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS2_OUT),
  .pad(`MP0_20),
  .pad_gz(`MP0_20_pad_y)
));
ap_MP0_20_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE)
));
ap_MP0_20_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_20_PINCTRL_0_IE),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_20),
  .pad(`MP0_20),
  .default_value(`default_value)));
ap_MP0_20_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_20_OUTFUNC_SEL),
  .gpioouten(`MP0_20_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`MP0_20_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`MP0_20),
  .pad_gz(`MP0_20_pad_y)
));
ap_MP0_20_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_20)
));
ap_MP0_20_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE)
));
ap_MP0_20_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_20_PINCTRL_0_IE),
  .outen(`MP0_20_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_20_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_20),
  .pad(`MP0_20),
  .default_value(`default_value)));
ap_MP0_20_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_20_PULLEN),
  .pullsel(`MP0_20_PULLSEL),
  .pad_pullup(`MP0_20)
));
ap_MP0_20_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .pullsel(`MP0_20_PULLSEL)
));
ap_MP0_20_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_20_PULLEN),
  .pullsel(`MP0_20_PULLSEL),
  .pad_pd(`MP0_20)
));
ap_MP0_20_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_20),
  .pullen(`MP0_20_PULLEN),
  .pullsel(`MP0_20_PULLSEL)
));
ap_MP0_21_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`MP0_21),
  .pad_gz(`MP0_21_pad_y)
));
ap_MP0_21_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE)
));
ap_MP0_21_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_21_PINCTRL_0_IE),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_21),
  .pad(`MP0_21),
  .default_value(`default_value)));
ap_MP0_21_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`MP0_21),
  .pad_gz(`MP0_21_pad_y)
));
ap_MP0_21_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE)
));
ap_MP0_21_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_21_PINCTRL_0_IE),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_21),
  .pad(`MP0_21),
  .default_value(`default_value)));
ap_MP0_21_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS3_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS3_OUT),
  .pad(`MP0_21),
  .pad_gz(`MP0_21_pad_y)
));
ap_MP0_21_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE)
));
ap_MP0_21_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_21_PINCTRL_0_IE),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_21),
  .pad(`MP0_21),
  .default_value(`default_value)));
ap_MP0_21_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_21_OUTFUNC_SEL),
  .gpioouten(`MP0_21_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`MP0_21_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`MP0_21),
  .pad_gz(`MP0_21_pad_y)
));
ap_MP0_21_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_21)
));
ap_MP0_21_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE)
));
ap_MP0_21_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_21_PINCTRL_0_IE),
  .outen(`MP0_21_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_21_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_21),
  .pad(`MP0_21),
  .default_value(`default_value)));
ap_MP0_21_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_21_PULLEN),
  .pullsel(`MP0_21_PULLSEL),
  .pad_pullup(`MP0_21)
));
ap_MP0_21_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .pullsel(`MP0_21_PULLSEL)
));
ap_MP0_21_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_21_PULLEN),
  .pullsel(`MP0_21_PULLSEL),
  .pad_pd(`MP0_21)
));
ap_MP0_21_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_21),
  .pullen(`MP0_21_PULLEN),
  .pullsel(`MP0_21_PULLSEL)
));
ap_MP0_22_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP0_22),
  .pad_gz(`MP0_22_pad_y)
));
ap_MP0_22_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_22),
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE)
));
ap_MP0_22_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_22_PINCTRL_0_IE),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_22),
  .pad(`MP0_22),
  .default_value(`default_value)));
ap_MP0_22_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`MP0_22),
  .pad_gz(`MP0_22_pad_y)
));
ap_MP0_22_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_22),
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE)
));
ap_MP0_22_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_22_PINCTRL_0_IE),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_22),
  .pad(`MP0_22),
  .default_value(`default_value)));
ap_MP0_22_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_22_OUTFUNC_SEL),
  .gpioouten(`MP0_22_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`MP0_22_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`MP0_22),
  .pad_gz(`MP0_22_pad_y)
));
ap_MP0_22_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_22)
));
ap_MP0_22_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_22),
  .pullen(`MP0_22_PULLEN),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE)
));
ap_MP0_22_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_22_PINCTRL_0_IE),
  .outen(`MP0_22_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_22_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_22),
  .pad(`MP0_22),
  .default_value(`default_value)));
ap_MP0_22_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_22_PULLEN),
  .pullsel(`MP0_22_PULLSEL),
  .pad_pullup(`MP0_22)
));
ap_MP0_22_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_22),
  .pullen(`MP0_22_PULLEN),
  .pullsel(`MP0_22_PULLSEL)
));
ap_MP0_22_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_22_PULLEN),
  .pullsel(`MP0_22_PULLSEL),
  .pad_pd(`MP0_22)
));
ap_MP0_22_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_22),
  .pullen(`MP0_22_PULLEN),
  .pullsel(`MP0_22_PULLSEL)
));
ap_MP0_23_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_23_OUTFUNC_SEL),
  .gpioouten(`MP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP0_23_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP0_23)
));
ap_MP0_23_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_23_OUTFUNC_SEL),
  .gpioouten(`MP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP0_23_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP0_23),
  .pad_gz(`MP0_23_pad_y)
));
ap_MP0_23_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_23_PULLEN),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_23)
));
ap_MP0_23_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_23),
  .pullen(`MP0_23_PULLEN),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE)
));
ap_MP0_23_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_23_PINCTRL_0_IE),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_23),
  .pad(`MP0_23),
  .default_value(`default_value)));
ap_MP0_23_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_23_OUTFUNC_SEL),
  .gpioouten(`MP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`MP0_23_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`MP0_23)
));
ap_MP0_23_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_23_OUTFUNC_SEL),
  .gpioouten(`MP0_23_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`MP0_23_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`MP0_23),
  .pad_gz(`MP0_23_pad_y)
));
ap_MP0_23_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_23_PULLEN),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_23)
));
ap_MP0_23_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_23),
  .pullen(`MP0_23_PULLEN),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE)
));
ap_MP0_23_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_23_PINCTRL_0_IE),
  .outen(`MP0_23_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_23_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_23),
  .pad(`MP0_23),
  .default_value(`default_value)));
ap_MP0_23_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_23_PULLEN),
  .pullsel(`MP0_23_PULLSEL),
  .pad_pullup(`MP0_23)
));
ap_MP0_23_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_23),
  .pullen(`MP0_23_PULLEN),
  .pullsel(`MP0_23_PULLSEL)
));
ap_MP0_23_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_23_PULLEN),
  .pullsel(`MP0_23_PULLSEL),
  .pad_pd(`MP0_23)
));
ap_MP0_23_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_23),
  .pullen(`MP0_23_PULLEN),
  .pullsel(`MP0_23_PULLSEL)
));
ap_MP0_24_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE)
));
ap_MP0_24_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_24_PINCTRL_0_IE),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_24),
  .pad(`MP0_24),
  .default_value(`default_value)));
ap_MP0_24_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_24_OUTFUNC_SEL),
  .gpioouten(`MP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`MP0_24_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_24_OUTFUNC_SEL),
  .gpioouten(`MP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`UART0TX_OE),
  .od(`MP0_24_PINCTRL_0_OD),
  .func_out(`UART0TX_OUT),
  .pad(`MP0_24),
  .pad_gz(`MP0_24_pad_y)
));
ap_MP0_24_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE)
));
ap_MP0_24_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_24_PINCTRL_0_IE),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_24),
  .pad(`MP0_24),
  .default_value(`default_value)));
ap_MP0_24_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE)
));
ap_MP0_24_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_24_PINCTRL_0_IE),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_24),
  .pad(`MP0_24),
  .default_value(`default_value)));
ap_MP0_24_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_24_OUTFUNC_SEL),
  .gpioouten(`MP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`MP0_24_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_24_OUTFUNC_SEL),
  .gpioouten(`MP0_24_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SDA_OE),
  .od(`MP0_24_PINCTRL_0_OD),
  .func_out(`I2C0SDA_OUT),
  .pad(`MP0_24),
  .pad_gz(`MP0_24_pad_y)
));
ap_MP0_24_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_24)
));
ap_MP0_24_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE)
));
ap_MP0_24_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_24_PINCTRL_0_IE),
  .outen(`MP0_24_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_24_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_24),
  .pad(`MP0_24),
  .default_value(`default_value)));
ap_MP0_24_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_24_PULLEN),
  .pullsel(`MP0_24_PULLSEL),
  .pad_pullup(`MP0_24)
));
ap_MP0_24_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .pullsel(`MP0_24_PULLSEL)
));
ap_MP0_24_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_24_PULLEN),
  .pullsel(`MP0_24_PULLSEL),
  .pad_pd(`MP0_24)
));
ap_MP0_24_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_24),
  .pullen(`MP0_24_PULLEN),
  .pullsel(`MP0_24_PULLSEL)
));
ap_MP0_25_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE)
));
ap_MP0_25_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_25_PINCTRL_0_IE),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_25),
  .pad(`MP0_25),
  .default_value(`default_value)));
ap_MP0_25_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_25_OUTFUNC_SEL),
  .gpioouten(`MP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`MP0_25_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_25_OUTFUNC_SEL),
  .gpioouten(`MP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`UART0RX_OE),
  .od(`MP0_25_PINCTRL_0_OD),
  .func_out(`UART0RX_OUT),
  .pad(`MP0_25),
  .pad_gz(`MP0_25_pad_y)
));
ap_MP0_25_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE)
));
ap_MP0_25_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_25_PINCTRL_0_IE),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_25),
  .pad(`MP0_25),
  .default_value(`default_value)));
ap_MP0_25_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE)
));
ap_MP0_25_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_25_PINCTRL_0_IE),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_25),
  .pad(`MP0_25),
  .default_value(`default_value)));
ap_MP0_25_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_25_OUTFUNC_SEL),
  .gpioouten(`MP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`MP0_25_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_25_OUTFUNC_SEL),
  .gpioouten(`MP0_25_GPIO_OUTPUT_ENABLE),
  .oe(`I2C0SCL_OE),
  .od(`MP0_25_PINCTRL_0_OD),
  .func_out(`I2C0SCL_OUT),
  .pad(`MP0_25),
  .pad_gz(`MP0_25_pad_y)
));
ap_MP0_25_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_25)
));
ap_MP0_25_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE)
));
ap_MP0_25_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_25_PINCTRL_0_IE),
  .outen(`MP0_25_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_25_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_25),
  .pad(`MP0_25),
  .default_value(`default_value)));
ap_MP0_25_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_25_PULLEN),
  .pullsel(`MP0_25_PULLSEL),
  .pad_pullup(`MP0_25)
));
ap_MP0_25_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .pullsel(`MP0_25_PULLSEL)
));
ap_MP0_25_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_25_PULLEN),
  .pullsel(`MP0_25_PULLSEL),
  .pad_pd(`MP0_25)
));
ap_MP0_25_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_25),
  .pullen(`MP0_25_PULLEN),
  .pullsel(`MP0_25_PULLSEL)
));
ap_MP0_26_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4TX_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`LIN4TX_OUT),
  .pad(`MP0_26),
  .pad_gz(`MP0_26_pad_y)
));
ap_MP0_26_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE)
));
ap_MP0_26_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_26_PINCTRL_0_IE),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_26),
  .pad(`MP0_26),
  .default_value(`default_value)));
ap_MP0_26_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`MP0_26),
  .pad_gz(`MP0_26_pad_y)
));
ap_MP0_26_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE)
));
ap_MP0_26_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_26_PINCTRL_0_IE),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_26),
  .pad(`MP0_26),
  .default_value(`default_value)));
ap_MP0_26_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE)
));
ap_MP0_26_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_26_PINCTRL_0_IE),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_26),
  .pad(`MP0_26),
  .default_value(`default_value)));
ap_MP0_26_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_26_OUTFUNC_SEL),
  .gpioouten(`MP0_26_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SDA_OE),
  .od(`MP0_26_PINCTRL_0_OD),
  .func_out(`I2C1SDA_OUT),
  .pad(`MP0_26),
  .pad_gz(`MP0_26_pad_y)
));
ap_MP0_26_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_26)
));
ap_MP0_26_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE)
));
ap_MP0_26_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_26_PINCTRL_0_IE),
  .outen(`MP0_26_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_26_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_26),
  .pad(`MP0_26),
  .default_value(`default_value)));
ap_MP0_26_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_26_PULLEN),
  .pullsel(`MP0_26_PULLSEL),
  .pad_pullup(`MP0_26)
));
ap_MP0_26_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .pullsel(`MP0_26_PULLSEL)
));
ap_MP0_26_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_26_PULLEN),
  .pullsel(`MP0_26_PULLSEL),
  .pad_pd(`MP0_26)
));
ap_MP0_26_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_26),
  .pullen(`MP0_26_PULLEN),
  .pullsel(`MP0_26_PULLSEL)
));
ap_MP0_27_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`LIN4RX_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`LIN4RX_OUT),
  .pad(`MP0_27),
  .pad_gz(`MP0_27_pad_y)
));
ap_MP0_27_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE)
));
ap_MP0_27_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_27_PINCTRL_0_IE),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_27),
  .pad(`MP0_27),
  .default_value(`default_value)));
ap_MP0_27_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`MP0_27),
  .pad_gz(`MP0_27_pad_y)
));
ap_MP0_27_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE)
));
ap_MP0_27_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_27_PINCTRL_0_IE),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_27),
  .pad(`MP0_27),
  .default_value(`default_value)));
ap_MP0_27_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE)
));
ap_MP0_27_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_27_PINCTRL_0_IE),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_27),
  .pad(`MP0_27),
  .default_value(`default_value)));
ap_MP0_27_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_27_OUTFUNC_SEL),
  .gpioouten(`MP0_27_GPIO_OUTPUT_ENABLE),
  .oe(`I2C1SCL_OE),
  .od(`MP0_27_PINCTRL_0_OD),
  .func_out(`I2C1SCL_OUT),
  .pad(`MP0_27),
  .pad_gz(`MP0_27_pad_y)
));
ap_MP0_27_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_27)
));
ap_MP0_27_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE)
));
ap_MP0_27_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_27_PINCTRL_0_IE),
  .outen(`MP0_27_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_27_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_27),
  .pad(`MP0_27),
  .default_value(`default_value)));
ap_MP0_27_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_27_PULLEN),
  .pullsel(`MP0_27_PULLSEL),
  .pad_pullup(`MP0_27)
));
ap_MP0_27_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .pullsel(`MP0_27_PULLSEL)
));
ap_MP0_27_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_27_PULLEN),
  .pullsel(`MP0_27_PULLSEL),
  .pad_pd(`MP0_27)
));
ap_MP0_27_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_27),
  .pullen(`MP0_27_PULLEN),
  .pullsel(`MP0_27_PULLSEL)
));
ap_MP0_28_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5TX_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`LIN5TX_OUT),
  .pad(`MP0_28),
  .pad_gz(`MP0_28_pad_y)
));
ap_MP0_28_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_28),
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE)
));
ap_MP0_28_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_28_PINCTRL_0_IE),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_28),
  .pad(`MP0_28),
  .default_value(`default_value)));
ap_MP0_28_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3TX_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`LIN3TX_OUT),
  .pad(`MP0_28),
  .pad_gz(`MP0_28_pad_y)
));
ap_MP0_28_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_28),
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE)
));
ap_MP0_28_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_28_PINCTRL_0_IE),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_28),
  .pad(`MP0_28),
  .default_value(`default_value)));
ap_MP0_28_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_28_OUTFUNC_SEL),
  .gpioouten(`MP0_28_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS11_OE),
  .od(`MP0_28_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS11_OUT),
  .pad(`MP0_28),
  .pad_gz(`MP0_28_pad_y)
));
ap_MP0_28_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_28)
));
ap_MP0_28_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_28),
  .pullen(`MP0_28_PULLEN),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE)
));
ap_MP0_28_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_28_PINCTRL_0_IE),
  .outen(`MP0_28_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_28_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_28),
  .pad(`MP0_28),
  .default_value(`default_value)));
ap_MP0_28_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_28_PULLEN),
  .pullsel(`MP0_28_PULLSEL),
  .pad_pullup(`MP0_28)
));
ap_MP0_28_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_28),
  .pullen(`MP0_28_PULLEN),
  .pullsel(`MP0_28_PULLSEL)
));
ap_MP0_28_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_28_PULLEN),
  .pullsel(`MP0_28_PULLSEL),
  .pad_pd(`MP0_28)
));
ap_MP0_28_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_28),
  .pullen(`MP0_28_PULLEN),
  .pullsel(`MP0_28_PULLSEL)
));
ap_MP0_29_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_29_OUTFUNC_SEL),
  .gpioouten(`MP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`MP0_29_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`MP0_29)
));
ap_MP0_29_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_29_OUTFUNC_SEL),
  .gpioouten(`MP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN5RX_OE),
  .od(`MP0_29_PINCTRL_0_OD),
  .func_out(`LIN5RX_OUT),
  .pad(`MP0_29),
  .pad_gz(`MP0_29_pad_y)
));
ap_MP0_29_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_29_PULLEN),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_29)
));
ap_MP0_29_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_29),
  .pullen(`MP0_29_PULLEN),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE)
));
ap_MP0_29_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_29_PINCTRL_0_IE),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_29_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_29),
  .pad(`MP0_29),
  .default_value(`default_value)));
ap_MP0_29_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_29_OUTFUNC_SEL),
  .gpioouten(`MP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`MP0_29_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`MP0_29)
));
ap_MP0_29_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_29_OUTFUNC_SEL),
  .gpioouten(`MP0_29_GPIO_OUTPUT_ENABLE),
  .oe(`LIN3RX_OE),
  .od(`MP0_29_PINCTRL_0_OD),
  .func_out(`LIN3RX_OUT),
  .pad(`MP0_29),
  .pad_gz(`MP0_29_pad_y)
));
ap_MP0_29_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_29_PULLEN),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_29)
));
ap_MP0_29_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_29),
  .pullen(`MP0_29_PULLEN),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE)
));
ap_MP0_29_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_29_PINCTRL_0_IE),
  .outen(`MP0_29_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_29_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_29),
  .pad(`MP0_29),
  .default_value(`default_value)));
ap_MP0_29_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_29_PULLEN),
  .pullsel(`MP0_29_PULLSEL),
  .pad_pullup(`MP0_29)
));
ap_MP0_29_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_29),
  .pullen(`MP0_29_PULLEN),
  .pullsel(`MP0_29_PULLSEL)
));
ap_MP0_29_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_29_PULLEN),
  .pullsel(`MP0_29_PULLSEL),
  .pad_pd(`MP0_29)
));
ap_MP0_29_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_29),
  .pullen(`MP0_29_PULLEN),
  .pullsel(`MP0_29_PULLSEL)
));
ap_MP0_30_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6TX_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`LIN6TX_OUT),
  .pad(`MP0_30),
  .pad_gz(`MP0_30_pad_y)
));
ap_MP0_30_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE)
));
ap_MP0_30_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_30_PINCTRL_0_IE),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_30),
  .pad(`MP0_30),
  .default_value(`default_value)));
ap_MP0_30_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS4_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`SPI6CS4_OUT),
  .pad(`MP0_30),
  .pad_gz(`MP0_30_pad_y)
));
ap_MP0_30_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE)
));
ap_MP0_30_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_30_PINCTRL_0_IE),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_30),
  .pad(`MP0_30),
  .default_value(`default_value)));
ap_MP0_30_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`MP0_30),
  .pad_gz(`MP0_30_pad_y)
));
ap_MP0_30_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE)
));
ap_MP0_30_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_30_PINCTRL_0_IE),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_30),
  .pad(`MP0_30),
  .default_value(`default_value)));
ap_MP0_30_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_30_OUTFUNC_SEL),
  .gpioouten(`MP0_30_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SDA_OE),
  .od(`MP0_30_PINCTRL_0_OD),
  .func_out(`I2C2SDA_OUT),
  .pad(`MP0_30),
  .pad_gz(`MP0_30_pad_y)
));
ap_MP0_30_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_30)
));
ap_MP0_30_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE)
));
ap_MP0_30_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_30_PINCTRL_0_IE),
  .outen(`MP0_30_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_30_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_30),
  .pad(`MP0_30),
  .default_value(`default_value)));
ap_MP0_30_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_30_PULLEN),
  .pullsel(`MP0_30_PULLSEL),
  .pad_pullup(`MP0_30)
));
ap_MP0_30_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .pullsel(`MP0_30_PULLSEL)
));
ap_MP0_30_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_30_PULLEN),
  .pullsel(`MP0_30_PULLSEL),
  .pad_pd(`MP0_30)
));
ap_MP0_30_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_30),
  .pullen(`MP0_30_PULLEN),
  .pullsel(`MP0_30_PULLSEL)
));
ap_MP0_31_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`LIN6RX_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`LIN6RX_OUT),
  .pad(`MP0_31),
  .pad_gz(`MP0_31_pad_y)
));
ap_MP0_31_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE)
));
ap_MP0_31_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP0_31_PINCTRL_0_IE),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_31),
  .pad(`MP0_31),
  .default_value(`default_value)));
ap_MP0_31_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`SPI6CS5_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`SPI6CS5_OUT),
  .pad(`MP0_31),
  .pad_gz(`MP0_31_pad_y)
));
ap_MP0_31_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE)
));
ap_MP0_31_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP0_31_PINCTRL_0_IE),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_31),
  .pad(`MP0_31),
  .default_value(`default_value)));
ap_MP0_31_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`MP0_31),
  .pad_gz(`MP0_31_pad_y)
));
ap_MP0_31_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE)
));
ap_MP0_31_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP0_31_PINCTRL_0_IE),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_31),
  .pad(`MP0_31),
  .default_value(`default_value)));
ap_MP0_31_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP0_31_OUTFUNC_SEL),
  .gpioouten(`MP0_31_GPIO_OUTPUT_ENABLE),
  .oe(`I2C2SCL_OE),
  .od(`MP0_31_PINCTRL_0_OD),
  .func_out(`I2C2SCL_OUT),
  .pad(`MP0_31),
  .pad_gz(`MP0_31_pad_y)
));
ap_MP0_31_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .pad(`MP0_31)
));
ap_MP0_31_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE)
));
ap_MP0_31_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP0_31_PINCTRL_0_IE),
  .outen(`MP0_31_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP0_31_INFUNC_EN),
  .in_concat(`input_func_concat_MP0_31),
  .pad(`MP0_31),
  .default_value(`default_value)));
ap_MP0_31_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP0_31_PULLEN),
  .pullsel(`MP0_31_PULLSEL),
  .pad_pullup(`MP0_31)
));
ap_MP0_31_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .pullsel(`MP0_31_PULLSEL)
));
ap_MP0_31_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP0_31_PULLEN),
  .pullsel(`MP0_31_PULLSEL),
  .pad_pd(`MP0_31)
));
ap_MP0_31_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP0_31),
  .pullen(`MP0_31_PULLEN),
  .pullsel(`MP0_31_PULLSEL)
));
ap_MP1_0_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7TX_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`LIN7TX_OUT),
  .pad(`MP1_0),
  .pad_gz(`MP1_0_pad_y)
));
ap_MP1_0_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE)
));
ap_MP1_0_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_0_PINCTRL_0_IE),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_0),
  .pad(`MP1_0),
  .default_value(`default_value)));
ap_MP1_0_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS4_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`SPI7CS4_OUT),
  .pad(`MP1_0),
  .pad_gz(`MP1_0_pad_y)
));
ap_MP1_0_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE)
));
ap_MP1_0_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_0_PINCTRL_0_IE),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_0),
  .pad(`MP1_0),
  .default_value(`default_value)));
ap_MP1_0_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`MP1_0),
  .pad_gz(`MP1_0_pad_y)
));
ap_MP1_0_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE)
));
ap_MP1_0_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP1_0_PINCTRL_0_IE),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_0),
  .pad(`MP1_0),
  .default_value(`default_value)));
ap_MP1_0_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_0_OUTFUNC_SEL),
  .gpioouten(`MP1_0_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SDA_OE),
  .od(`MP1_0_PINCTRL_0_OD),
  .func_out(`I2C3SDA_OUT),
  .pad(`MP1_0),
  .pad_gz(`MP1_0_pad_y)
));
ap_MP1_0_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_0)
));
ap_MP1_0_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE)
));
ap_MP1_0_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP1_0_PINCTRL_0_IE),
  .outen(`MP1_0_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_0_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_0),
  .pad(`MP1_0),
  .default_value(`default_value)));
ap_MP1_0_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_0_PULLEN),
  .pullsel(`MP1_0_PULLSEL),
  .pad_pullup(`MP1_0)
));
ap_MP1_0_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .pullsel(`MP1_0_PULLSEL)
));
ap_MP1_0_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_0_PULLEN),
  .pullsel(`MP1_0_PULLSEL),
  .pad_pd(`MP1_0)
));
ap_MP1_0_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_0),
  .pullen(`MP1_0_PULLEN),
  .pullsel(`MP1_0_PULLSEL)
));
ap_MP1_1_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`LIN7RX_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`LIN7RX_OUT),
  .pad(`MP1_1),
  .pad_gz(`MP1_1_pad_y)
));
ap_MP1_1_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE)
));
ap_MP1_1_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_1_PINCTRL_0_IE),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_1),
  .pad(`MP1_1),
  .default_value(`default_value)));
ap_MP1_1_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`SPI7CS5_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`SPI7CS5_OUT),
  .pad(`MP1_1),
  .pad_gz(`MP1_1_pad_y)
));
ap_MP1_1_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE)
));
ap_MP1_1_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_1_PINCTRL_0_IE),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_1),
  .pad(`MP1_1),
  .default_value(`default_value)));
ap_MP1_1_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS8_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS8_OUT),
  .pad(`MP1_1),
  .pad_gz(`MP1_1_pad_y)
));
ap_MP1_1_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE)
));
ap_MP1_1_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP1_1_PINCTRL_0_IE),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_1),
  .pad(`MP1_1),
  .default_value(`default_value)));
ap_MP1_1_FUNCSEL_4_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_4_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_1_OUTFUNC_SEL),
  .gpioouten(`MP1_1_GPIO_OUTPUT_ENABLE),
  .oe(`I2C3SCL_OE),
  .od(`MP1_1_PINCTRL_0_OD),
  .func_out(`I2C3SCL_OUT),
  .pad(`MP1_1),
  .pad_gz(`MP1_1_pad_y)
));
ap_MP1_1_FUNCSEL_4_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_1)
));
ap_MP1_1_FUNCSEL_4_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE)
));
ap_MP1_1_FUNCSEL_4_input_chk : assert property(iomux_input_path(
  .ie(`MP1_1_PINCTRL_0_IE),
  .outen(`MP1_1_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_1_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_1),
  .pad(`MP1_1),
  .default_value(`default_value)));
ap_MP1_1_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_1_PULLEN),
  .pullsel(`MP1_1_PULLSEL),
  .pad_pullup(`MP1_1)
));
ap_MP1_1_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .pullsel(`MP1_1_PULLSEL)
));
ap_MP1_1_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_1_PULLEN),
  .pullsel(`MP1_1_PULLSEL),
  .pad_pd(`MP1_1)
));
ap_MP1_1_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_1),
  .pullen(`MP1_1_PULLEN),
  .pullsel(`MP1_1_PULLSEL)
));
ap_MP1_2_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`UART1TX_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`UART1TX_OUT),
  .pad(`MP1_2),
  .pad_gz(`MP1_2_pad_y)
));
ap_MP1_2_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_2),
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE)
));
ap_MP1_2_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_2_PINCTRL_0_IE),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_2),
  .pad(`MP1_2),
  .default_value(`default_value)));
ap_MP1_2_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP1_2),
  .pad_gz(`MP1_2_pad_y)
));
ap_MP1_2_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_2),
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE)
));
ap_MP1_2_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_2_PINCTRL_0_IE),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_2),
  .pad(`MP1_2),
  .default_value(`default_value)));
ap_MP1_2_FUNCSEL_3_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_3_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_2_OUTFUNC_SEL),
  .gpioouten(`MP1_2_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS9_OE),
  .od(`MP1_2_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS9_OUT),
  .pad(`MP1_2),
  .pad_gz(`MP1_2_pad_y)
));
ap_MP1_2_FUNCSEL_3_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_2)
));
ap_MP1_2_FUNCSEL_3_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_2),
  .pullen(`MP1_2_PULLEN),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE)
));
ap_MP1_2_FUNCSEL_3_input_chk : assert property(iomux_input_path(
  .ie(`MP1_2_PINCTRL_0_IE),
  .outen(`MP1_2_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_2_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_2),
  .pad(`MP1_2),
  .default_value(`default_value)));
ap_MP1_2_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_2_PULLEN),
  .pullsel(`MP1_2_PULLSEL),
  .pad_pullup(`MP1_2)
));
ap_MP1_2_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_2),
  .pullen(`MP1_2_PULLEN),
  .pullsel(`MP1_2_PULLSEL)
));
ap_MP1_2_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_2_PULLEN),
  .pullsel(`MP1_2_PULLSEL),
  .pad_pd(`MP1_2)
));
ap_MP1_2_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_2),
  .pullen(`MP1_2_PULLEN),
  .pullsel(`MP1_2_PULLSEL)
));
ap_MP1_3_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_3_OUTFUNC_SEL),
  .gpioouten(`MP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`MP1_3_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`MP1_3)
));
ap_MP1_3_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_3_OUTFUNC_SEL),
  .gpioouten(`MP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`UART1RX_OE),
  .od(`MP1_3_PINCTRL_0_OD),
  .func_out(`UART1RX_OUT),
  .pad(`MP1_3),
  .pad_gz(`MP1_3_pad_y)
));
ap_MP1_3_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_3_PULLEN),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_3)
));
ap_MP1_3_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_3),
  .pullen(`MP1_3_PULLEN),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE)
));
ap_MP1_3_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_3_PINCTRL_0_IE),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_3),
  .pad(`MP1_3),
  .default_value(`default_value)));
ap_MP1_3_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_3_OUTFUNC_SEL),
  .gpioouten(`MP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP1_3_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP1_3)
));
ap_MP1_3_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_3_OUTFUNC_SEL),
  .gpioouten(`MP1_3_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP1_3_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP1_3),
  .pad_gz(`MP1_3_pad_y)
));
ap_MP1_3_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_3_PULLEN),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_3)
));
ap_MP1_3_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_3),
  .pullen(`MP1_3_PULLEN),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE)
));
ap_MP1_3_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_3_PINCTRL_0_IE),
  .outen(`MP1_3_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_3_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_3),
  .pad(`MP1_3),
  .default_value(`default_value)));
ap_MP1_3_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_3_PULLEN),
  .pullsel(`MP1_3_PULLSEL),
  .pad_pullup(`MP1_3)
));
ap_MP1_3_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_3),
  .pullen(`MP1_3_PULLEN),
  .pullsel(`MP1_3_PULLSEL)
));
ap_MP1_3_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_3_PULLEN),
  .pullsel(`MP1_3_PULLSEL),
  .pad_pd(`MP1_3)
));
ap_MP1_3_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_3),
  .pullen(`MP1_3_PULLEN),
  .pullsel(`MP1_3_PULLSEL)
));
ap_MP1_4_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_4_OUTFUNC_SEL),
  .gpioouten(`MP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`MP1_4_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`MP1_4)
));
ap_MP1_4_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_4_OUTFUNC_SEL),
  .gpioouten(`MP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`SENT0TXRX_OE),
  .od(`MP1_4_PINCTRL_0_OD),
  .func_out(`SENT0TXRX_OUT),
  .pad(`MP1_4),
  .pad_gz(`MP1_4_pad_y)
));
ap_MP1_4_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_4_PULLEN),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_4)
));
ap_MP1_4_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_4),
  .pullen(`MP1_4_PULLEN),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE)
));
ap_MP1_4_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_4_PINCTRL_0_IE),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_4),
  .pad(`MP1_4),
  .default_value(`default_value)));
ap_MP1_4_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_4_OUTFUNC_SEL),
  .gpioouten(`MP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP1_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP1_4)
));
ap_MP1_4_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_4_OUTFUNC_SEL),
  .gpioouten(`MP1_4_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS4_OE),
  .od(`MP1_4_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS4_OUT),
  .pad(`MP1_4),
  .pad_gz(`MP1_4_pad_y)
));
ap_MP1_4_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_4_PULLEN),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_4)
));
ap_MP1_4_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_4),
  .pullen(`MP1_4_PULLEN),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE)
));
ap_MP1_4_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_4_PINCTRL_0_IE),
  .outen(`MP1_4_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_4_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_4),
  .pad(`MP1_4),
  .default_value(`default_value)));
ap_MP1_4_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_4_PULLEN),
  .pullsel(`MP1_4_PULLSEL),
  .pad_pullup(`MP1_4)
));
ap_MP1_4_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_4),
  .pullen(`MP1_4_PULLEN),
  .pullsel(`MP1_4_PULLSEL)
));
ap_MP1_4_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_4_PULLEN),
  .pullsel(`MP1_4_PULLSEL),
  .pad_pd(`MP1_4)
));
ap_MP1_4_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_4),
  .pullen(`MP1_4_PULLEN),
  .pullsel(`MP1_4_PULLSEL)
));
ap_MP1_5_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_5_OUTFUNC_SEL),
  .gpioouten(`MP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`MP1_5_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`MP1_5)
));
ap_MP1_5_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_5_OUTFUNC_SEL),
  .gpioouten(`MP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`SENT1TXRX_OE),
  .od(`MP1_5_PINCTRL_0_OD),
  .func_out(`SENT1TXRX_OUT),
  .pad(`MP1_5),
  .pad_gz(`MP1_5_pad_y)
));
ap_MP1_5_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_5_PULLEN),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_5)
));
ap_MP1_5_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_5),
  .pullen(`MP1_5_PULLEN),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE)
));
ap_MP1_5_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_5_PINCTRL_0_IE),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_5),
  .pad(`MP1_5),
  .default_value(`default_value)));
ap_MP1_5_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_5_OUTFUNC_SEL),
  .gpioouten(`MP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP1_5_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP1_5)
));
ap_MP1_5_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_5_OUTFUNC_SEL),
  .gpioouten(`MP1_5_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS5_OE),
  .od(`MP1_5_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS5_OUT),
  .pad(`MP1_5),
  .pad_gz(`MP1_5_pad_y)
));
ap_MP1_5_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_5_PULLEN),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_5)
));
ap_MP1_5_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_5),
  .pullen(`MP1_5_PULLEN),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE)
));
ap_MP1_5_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_5_PINCTRL_0_IE),
  .outen(`MP1_5_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_5_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_5),
  .pad(`MP1_5),
  .default_value(`default_value)));
ap_MP1_5_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_5_PULLEN),
  .pullsel(`MP1_5_PULLSEL),
  .pad_pullup(`MP1_5)
));
ap_MP1_5_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_5),
  .pullen(`MP1_5_PULLEN),
  .pullsel(`MP1_5_PULLSEL)
));
ap_MP1_5_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_5_PULLEN),
  .pullsel(`MP1_5_PULLSEL),
  .pad_pd(`MP1_5)
));
ap_MP1_5_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_5),
  .pullen(`MP1_5_PULLEN),
  .pullsel(`MP1_5_PULLSEL)
));
ap_MP1_6_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_6_OUTFUNC_SEL),
  .gpioouten(`MP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`MP1_6_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`MP1_6)
));
ap_MP1_6_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_6_OUTFUNC_SEL),
  .gpioouten(`MP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`SENT2TXRX_OE),
  .od(`MP1_6_PINCTRL_0_OD),
  .func_out(`SENT2TXRX_OUT),
  .pad(`MP1_6),
  .pad_gz(`MP1_6_pad_y)
));
ap_MP1_6_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_6_PULLEN),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_6)
));
ap_MP1_6_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_6),
  .pullen(`MP1_6_PULLEN),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE)
));
ap_MP1_6_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_6_PINCTRL_0_IE),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_6),
  .pad(`MP1_6),
  .default_value(`default_value)));
ap_MP1_6_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_6_OUTFUNC_SEL),
  .gpioouten(`MP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP1_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP1_6)
));
ap_MP1_6_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_6_OUTFUNC_SEL),
  .gpioouten(`MP1_6_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS6_OE),
  .od(`MP1_6_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS6_OUT),
  .pad(`MP1_6),
  .pad_gz(`MP1_6_pad_y)
));
ap_MP1_6_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_6_PULLEN),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_6)
));
ap_MP1_6_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_6),
  .pullen(`MP1_6_PULLEN),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE)
));
ap_MP1_6_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_6_PINCTRL_0_IE),
  .outen(`MP1_6_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_6_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_6),
  .pad(`MP1_6),
  .default_value(`default_value)));
ap_MP1_6_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_6_PULLEN),
  .pullsel(`MP1_6_PULLSEL),
  .pad_pullup(`MP1_6)
));
ap_MP1_6_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_6),
  .pullen(`MP1_6_PULLEN),
  .pullsel(`MP1_6_PULLSEL)
));
ap_MP1_6_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_6_PULLEN),
  .pullsel(`MP1_6_PULLSEL),
  .pad_pd(`MP1_6)
));
ap_MP1_6_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_6),
  .pullen(`MP1_6_PULLEN),
  .pullsel(`MP1_6_PULLSEL)
));
ap_MP1_7_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_7_OUTFUNC_SEL),
  .gpioouten(`MP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`MP1_7_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`MP1_7)
));
ap_MP1_7_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_7_OUTFUNC_SEL),
  .gpioouten(`MP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`SENT3TXRX_OE),
  .od(`MP1_7_PINCTRL_0_OD),
  .func_out(`SENT3TXRX_OUT),
  .pad(`MP1_7),
  .pad_gz(`MP1_7_pad_y)
));
ap_MP1_7_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_7_PULLEN),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_7)
));
ap_MP1_7_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_7),
  .pullen(`MP1_7_PULLEN),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE)
));
ap_MP1_7_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_7_PINCTRL_0_IE),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_7),
  .pad(`MP1_7),
  .default_value(`default_value)));
ap_MP1_7_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_7_OUTFUNC_SEL),
  .gpioouten(`MP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP1_7_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP1_7)
));
ap_MP1_7_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_7_OUTFUNC_SEL),
  .gpioouten(`MP1_7_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS7_OE),
  .od(`MP1_7_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS7_OUT),
  .pad(`MP1_7),
  .pad_gz(`MP1_7_pad_y)
));
ap_MP1_7_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_7_PULLEN),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_7)
));
ap_MP1_7_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_7),
  .pullen(`MP1_7_PULLEN),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE)
));
ap_MP1_7_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_7_PINCTRL_0_IE),
  .outen(`MP1_7_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_7_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_7),
  .pad(`MP1_7),
  .default_value(`default_value)));
ap_MP1_7_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_7_PULLEN),
  .pullsel(`MP1_7_PULLSEL),
  .pad_pullup(`MP1_7)
));
ap_MP1_7_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_7),
  .pullen(`MP1_7_PULLEN),
  .pullsel(`MP1_7_PULLSEL)
));
ap_MP1_7_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_7_PULLEN),
  .pullsel(`MP1_7_PULLSEL),
  .pad_pd(`MP1_7)
));
ap_MP1_7_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_7),
  .pullen(`MP1_7_PULLEN),
  .pullsel(`MP1_7_PULLSEL)
));
ap_MP1_8_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_8_OUTFUNC_SEL),
  .gpioouten(`MP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP1_8_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP1_8)
));
ap_MP1_8_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_8_OUTFUNC_SEL),
  .gpioouten(`MP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`SENT4TXRX_OE),
  .od(`MP1_8_PINCTRL_0_OD),
  .func_out(`SENT4TXRX_OUT),
  .pad(`MP1_8),
  .pad_gz(`MP1_8_pad_y)
));
ap_MP1_8_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_8_PULLEN),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_8)
));
ap_MP1_8_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_8),
  .pullen(`MP1_8_PULLEN),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE)
));
ap_MP1_8_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_8_PINCTRL_0_IE),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_8),
  .pad(`MP1_8),
  .default_value(`default_value)));
ap_MP1_8_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_8_OUTFUNC_SEL),
  .gpioouten(`MP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP1_8_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP1_8)
));
ap_MP1_8_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_8_OUTFUNC_SEL),
  .gpioouten(`MP1_8_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS8_OE),
  .od(`MP1_8_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS8_OUT),
  .pad(`MP1_8),
  .pad_gz(`MP1_8_pad_y)
));
ap_MP1_8_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_8_PULLEN),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_8)
));
ap_MP1_8_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_8),
  .pullen(`MP1_8_PULLEN),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE)
));
ap_MP1_8_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_8_PINCTRL_0_IE),
  .outen(`MP1_8_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_8_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_8),
  .pad(`MP1_8),
  .default_value(`default_value)));
ap_MP1_8_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_8_PULLEN),
  .pullsel(`MP1_8_PULLSEL),
  .pad_pullup(`MP1_8)
));
ap_MP1_8_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_8),
  .pullen(`MP1_8_PULLEN),
  .pullsel(`MP1_8_PULLSEL)
));
ap_MP1_8_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_8_PULLEN),
  .pullsel(`MP1_8_PULLSEL),
  .pad_pd(`MP1_8)
));
ap_MP1_8_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_8),
  .pullen(`MP1_8_PULLEN),
  .pullsel(`MP1_8_PULLSEL)
));
ap_MP1_9_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_9_OUTFUNC_SEL),
  .gpioouten(`MP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP1_9_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP1_9)
));
ap_MP1_9_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_9_OUTFUNC_SEL),
  .gpioouten(`MP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`SENT5TXRX_OE),
  .od(`MP1_9_PINCTRL_0_OD),
  .func_out(`SENT5TXRX_OUT),
  .pad(`MP1_9),
  .pad_gz(`MP1_9_pad_y)
));
ap_MP1_9_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_9_PULLEN),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_9)
));
ap_MP1_9_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_9),
  .pullen(`MP1_9_PULLEN),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE)
));
ap_MP1_9_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_9_PINCTRL_0_IE),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_9),
  .pad(`MP1_9),
  .default_value(`default_value)));
ap_MP1_9_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_9_OUTFUNC_SEL),
  .gpioouten(`MP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP1_9_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP1_9)
));
ap_MP1_9_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_9_OUTFUNC_SEL),
  .gpioouten(`MP1_9_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS9_OE),
  .od(`MP1_9_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS9_OUT),
  .pad(`MP1_9),
  .pad_gz(`MP1_9_pad_y)
));
ap_MP1_9_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_9_PULLEN),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_9)
));
ap_MP1_9_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_9),
  .pullen(`MP1_9_PULLEN),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE)
));
ap_MP1_9_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_9_PINCTRL_0_IE),
  .outen(`MP1_9_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_9_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_9),
  .pad(`MP1_9),
  .default_value(`default_value)));
ap_MP1_9_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_9_PULLEN),
  .pullsel(`MP1_9_PULLSEL),
  .pad_pullup(`MP1_9)
));
ap_MP1_9_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_9),
  .pullen(`MP1_9_PULLEN),
  .pullsel(`MP1_9_PULLSEL)
));
ap_MP1_9_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_9_PULLEN),
  .pullsel(`MP1_9_PULLSEL),
  .pad_pd(`MP1_9)
));
ap_MP1_9_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_9),
  .pullen(`MP1_9_PULLEN),
  .pullsel(`MP1_9_PULLSEL)
));
ap_MP1_10_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_10_OUTFUNC_SEL),
  .gpioouten(`MP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`MP1_10_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`MP1_10)
));
ap_MP1_10_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_10_OUTFUNC_SEL),
  .gpioouten(`MP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS4_OE),
  .od(`MP1_10_PINCTRL_0_OD),
  .func_out(`SPI5CS4_OUT),
  .pad(`MP1_10),
  .pad_gz(`MP1_10_pad_y)
));
ap_MP1_10_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_10_PULLEN),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_10)
));
ap_MP1_10_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_10),
  .pullen(`MP1_10_PULLEN),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE)
));
ap_MP1_10_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_10_PINCTRL_0_IE),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_10),
  .pad(`MP1_10),
  .default_value(`default_value)));
ap_MP1_10_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_10_OUTFUNC_SEL),
  .gpioouten(`MP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP1_10_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP1_10)
));
ap_MP1_10_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_10_OUTFUNC_SEL),
  .gpioouten(`MP1_10_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS10_OE),
  .od(`MP1_10_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS10_OUT),
  .pad(`MP1_10),
  .pad_gz(`MP1_10_pad_y)
));
ap_MP1_10_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_10_PULLEN),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_10)
));
ap_MP1_10_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_10),
  .pullen(`MP1_10_PULLEN),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE)
));
ap_MP1_10_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_10_PINCTRL_0_IE),
  .outen(`MP1_10_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_10_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_10),
  .pad(`MP1_10),
  .default_value(`default_value)));
ap_MP1_10_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_10_PULLEN),
  .pullsel(`MP1_10_PULLSEL),
  .pad_pullup(`MP1_10)
));
ap_MP1_10_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_10),
  .pullen(`MP1_10_PULLEN),
  .pullsel(`MP1_10_PULLSEL)
));
ap_MP1_10_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_10_PULLEN),
  .pullsel(`MP1_10_PULLSEL),
  .pad_pd(`MP1_10)
));
ap_MP1_10_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_10),
  .pullen(`MP1_10_PULLEN),
  .pullsel(`MP1_10_PULLSEL)
));
ap_MP1_11_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_11_OUTFUNC_SEL),
  .gpioouten(`MP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`MP1_11_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`MP1_11)
));
ap_MP1_11_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_11_OUTFUNC_SEL),
  .gpioouten(`MP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`SPI5CS5_OE),
  .od(`MP1_11_PINCTRL_0_OD),
  .func_out(`SPI5CS5_OUT),
  .pad(`MP1_11),
  .pad_gz(`MP1_11_pad_y)
));
ap_MP1_11_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_11_PULLEN),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_11)
));
ap_MP1_11_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_11),
  .pullen(`MP1_11_PULLEN),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE)
));
ap_MP1_11_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_11_PINCTRL_0_IE),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_11),
  .pad(`MP1_11),
  .default_value(`default_value)));
ap_MP1_11_FUNCSEL_2_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_11_OUTFUNC_SEL),
  .gpioouten(`MP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP1_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP1_11)
));
ap_MP1_11_FUNCSEL_2_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_11_OUTFUNC_SEL),
  .gpioouten(`MP1_11_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI1CS11_OE),
  .od(`MP1_11_PINCTRL_0_OD),
  .func_out(`MIBSPI1CS11_OUT),
  .pad(`MP1_11),
  .pad_gz(`MP1_11_pad_y)
));
ap_MP1_11_FUNCSEL_2_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_11_PULLEN),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_11)
));
ap_MP1_11_FUNCSEL_2_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_11),
  .pullen(`MP1_11_PULLEN),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE)
));
ap_MP1_11_FUNCSEL_2_input_chk : assert property(iomux_input_path(
  .ie(`MP1_11_PINCTRL_0_IE),
  .outen(`MP1_11_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_11_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_11),
  .pad(`MP1_11),
  .default_value(`default_value)));
ap_MP1_11_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_11_PULLEN),
  .pullsel(`MP1_11_PULLSEL),
  .pad_pullup(`MP1_11)
));
ap_MP1_11_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_11),
  .pullen(`MP1_11_PULLEN),
  .pullsel(`MP1_11_PULLSEL)
));
ap_MP1_11_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_11_PULLEN),
  .pullsel(`MP1_11_PULLSEL),
  .pad_pd(`MP1_11)
));
ap_MP1_11_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_11),
  .pullen(`MP1_11_PULLEN),
  .pullsel(`MP1_11_PULLSEL)
));
ap_MP1_12_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_12_OUTFUNC_SEL),
  .gpioouten(`MP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`MP1_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`MP1_12)
));
ap_MP1_12_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_12_OUTFUNC_SEL),
  .gpioouten(`MP1_12_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS4_OE),
  .od(`MP1_12_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS4_OUT),
  .pad(`MP1_12),
  .pad_gz(`MP1_12_pad_y)
));
ap_MP1_12_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_12_PULLEN),
  .outen(`MP1_12_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_12)
));
ap_MP1_12_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_12),
  .pullen(`MP1_12_PULLEN),
  .outen(`MP1_12_GPIO_OUTPUT_ENABLE)
));
ap_MP1_12_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_12_PINCTRL_0_IE),
  .outen(`MP1_12_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_12_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_12),
  .pad(`MP1_12),
  .default_value(`default_value)));
ap_MP1_12_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_12_PULLEN),
  .pullsel(`MP1_12_PULLSEL),
  .pad_pullup(`MP1_12)
));
ap_MP1_12_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_12),
  .pullen(`MP1_12_PULLEN),
  .pullsel(`MP1_12_PULLSEL)
));
ap_MP1_12_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_12_PULLEN),
  .pullsel(`MP1_12_PULLSEL),
  .pad_pd(`MP1_12)
));
ap_MP1_12_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_12),
  .pullen(`MP1_12_PULLEN),
  .pullsel(`MP1_12_PULLSEL)
));
ap_MP1_13_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_13_OUTFUNC_SEL),
  .gpioouten(`MP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`MP1_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`MP1_13)
));
ap_MP1_13_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_13_OUTFUNC_SEL),
  .gpioouten(`MP1_13_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS5_OE),
  .od(`MP1_13_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS5_OUT),
  .pad(`MP1_13),
  .pad_gz(`MP1_13_pad_y)
));
ap_MP1_13_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_13_PULLEN),
  .outen(`MP1_13_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_13)
));
ap_MP1_13_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_13),
  .pullen(`MP1_13_PULLEN),
  .outen(`MP1_13_GPIO_OUTPUT_ENABLE)
));
ap_MP1_13_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_13_PINCTRL_0_IE),
  .outen(`MP1_13_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_13_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_13),
  .pad(`MP1_13),
  .default_value(`default_value)));
ap_MP1_13_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_13_PULLEN),
  .pullsel(`MP1_13_PULLSEL),
  .pad_pullup(`MP1_13)
));
ap_MP1_13_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_13),
  .pullen(`MP1_13_PULLEN),
  .pullsel(`MP1_13_PULLSEL)
));
ap_MP1_13_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_13_PULLEN),
  .pullsel(`MP1_13_PULLSEL),
  .pad_pd(`MP1_13)
));
ap_MP1_13_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_13),
  .pullen(`MP1_13_PULLEN),
  .pullsel(`MP1_13_PULLSEL)
));
ap_MP1_14_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_14_OUTFUNC_SEL),
  .gpioouten(`MP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`MP1_14_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`MP1_14)
));
ap_MP1_14_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_14_OUTFUNC_SEL),
  .gpioouten(`MP1_14_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS6_OE),
  .od(`MP1_14_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS6_OUT),
  .pad(`MP1_14),
  .pad_gz(`MP1_14_pad_y)
));
ap_MP1_14_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_14_PULLEN),
  .outen(`MP1_14_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_14)
));
ap_MP1_14_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_14),
  .pullen(`MP1_14_PULLEN),
  .outen(`MP1_14_GPIO_OUTPUT_ENABLE)
));
ap_MP1_14_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_14_PINCTRL_0_IE),
  .outen(`MP1_14_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_14_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_14),
  .pad(`MP1_14),
  .default_value(`default_value)));
ap_MP1_14_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_14_PULLEN),
  .pullsel(`MP1_14_PULLSEL),
  .pad_pullup(`MP1_14)
));
ap_MP1_14_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_14),
  .pullen(`MP1_14_PULLEN),
  .pullsel(`MP1_14_PULLSEL)
));
ap_MP1_14_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_14_PULLEN),
  .pullsel(`MP1_14_PULLSEL),
  .pad_pd(`MP1_14)
));
ap_MP1_14_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_14),
  .pullen(`MP1_14_PULLEN),
  .pullsel(`MP1_14_PULLSEL)
));
ap_MP1_15_FUNCSEL_1_output_drive_chk : assert property(iomux_output_drive(
  .funcsel(`MP1_15_OUTFUNC_SEL),
  .gpioouten(`MP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`MP1_15_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`MP1_15)
));
ap_MP1_15_FUNCSEL_1_open_drain_chk : assert property(iomux_output_open_drain(
  .funcsel(`MP1_15_OUTFUNC_SEL),
  .gpioouten(`MP1_15_GPIO_OUTPUT_ENABLE),
  .oe(`MIBSPI0CS7_OE),
  .od(`MP1_15_PINCTRL_0_OD),
  .func_out(`MIBSPI0CS7_OUT),
  .pad(`MP1_15),
  .pad_gz(`MP1_15_pad_y)
));
ap_MP1_15_FUNCSEL_1_highz_cond_chk : assert property(iomux_highz_conditions(
  .pullen(`MP1_15_PULLEN),
  .outen(`MP1_15_GPIO_OUTPUT_ENABLE),
  .pad(`MP1_15)
));
ap_MP1_15_FUNCSEL_1_highz_rev_chk : assert property(iomux_highz_reverse(
  .pad(`MP1_15),
  .pullen(`MP1_15_PULLEN),
  .outen(`MP1_15_GPIO_OUTPUT_ENABLE)
));
ap_MP1_15_FUNCSEL_1_input_chk : assert property(iomux_input_path(
  .ie(`MP1_15_PINCTRL_0_IE),
  .outen(`MP1_15_GPIO_OUTPUT_ENABLE),
  .infunc_en(`MP1_15_INFUNC_EN),
  .in_concat(`input_func_concat_MP1_15),
  .pad(`MP1_15),
  .default_value(`default_value)));
ap_MP1_15_FUNCSEL_pull_up_chk : assert property(iomux_pull_up(
  .pullen(`MP1_15_PULLEN),
  .pullsel(`MP1_15_PULLSEL),
  .pad_pullup(`MP1_15)
));
ap_MP1_15_FUNCSEL_pull_up_reverse_chk : assert property(iomux_pull_up_reverse(
  .pad_pullup(`MP1_15),
  .pullen(`MP1_15_PULLEN),
  .pullsel(`MP1_15_PULLSEL)
));
ap_MP1_15_FUNCSEL_pull_down_chk : assert property(iomux_pull_down(
  .pullen(`MP1_15_PULLEN),
  .pullsel(`MP1_15_PULLSEL),
  .pad_pd(`MP1_15)
));
ap_MP1_15_FUNCSEL_pull_down_reverse_chk : assert property(iomux_pull_down_reverse(
  .pad_pd(`MP1_15),
  .pullen(`MP1_15_PULLEN),
  .pullsel(`MP1_15_PULLSEL)
));

endmodule

bind assertion_gen pinmux_wrapper bind_inst();
