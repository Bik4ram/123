//====================================================================
// Copyright (c) 2025 Texas Instruments, Inc.
// This is an unpublished work created in the year stated above.
// Texas Instruments owns all rights in and to this work and
// intends to maintain and protect it as an unpublished copyright.
// In the event of either inadvertent or deliberate publication,
// the above stated date shall be treated as the year of first
// publication. In the event of such publication, Texas Instruments
// intends to enforce its rights in the work under the copyright
// laws as a published work.
//====================================================================
//
// pinmux_wrapper.v
//
//    pinmux wrapper
//
//====================================================================
// Module Designer: Himanshi (h-himanshi@ti.com)
// Contact Info:    Texas Instruments
//                  DSP Systems /  Group
//                  12500 TI Blvd
//                  Dallas, Texas 75243
//                  (918)708-488241
//
//====================================================================
// Revision History:
//  1.0.0.0 15/1/2025 spec a0507242 first version
//
//====================================================================
// Generated by VeriPerl Compiler version 3.0.347
//    Build 2021.09.22.09.59.05
//
//====================================================================
`timescale 1 ps / 1 ps


module pinmux_wrapper (

  // dp0 async input from pad bus
  dp0_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp0 gpio out to buf bus
  dp0_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp0 gpio out enable bus
  dp0_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp0 pinmux data to gpio bus
  dp0_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp0 pinmux enable to gpio bus
  dp0_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp0 GP DATA IN out bus
  dp0_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp0 data out to pinmux bus
  dp0_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp0 pinmux muxsel out bus
  dp0_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp0 in function enable out bus
  dp0_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp0 analog mode select bus
  dp0_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp0 drive strength 0 bus
  dp0_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp0 drive strength 1 bus
  dp0_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp0 slew control bus
  dp0_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp0 schmitt trigger bus
  dp0_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp0 mode 0 bus
  dp0_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp0 mode 1 bus
  dp0_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp0 input enable bus
  dp0_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp0 direction bus
  dp0_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp0 pull enable bus
  dp0_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp0 pull type bus
  dp0_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp0 glitch filter debounce clock select bus
  dp0_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp0 glitch filter bypass bus
  dp0_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp0 PES enable bus
  dp0_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp0 PES input enable bus
  dp0_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp0 PES safe value bus
  dp0_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp0 LVDS enable control bus
  dp0_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp0 input termination enable bus
  dp0_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp1 async input from pad bus
  dp1_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp1 gpio out to buf bus
  dp1_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp1 gpio out enable bus
  dp1_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp1 pinmux data to gpio bus
  dp1_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp1 pinmux enable to gpio bus
  dp1_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp1 GP DATA IN out bus
  dp1_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp1 data out to pinmux bus
  dp1_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp1 pinmux muxsel out bus
  dp1_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp1 in function enable out bus
  dp1_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp1 analog mode select bus
  dp1_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp1 drive strength 0 bus
  dp1_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp1 drive strength 1 bus
  dp1_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp1 slew control bus
  dp1_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp1 schmitt trigger bus
  dp1_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp1 mode 0 bus
  dp1_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp1 mode 1 bus
  dp1_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp1 input enable bus
  dp1_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp1 direction bus
  dp1_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp1 pull enable bus
  dp1_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp1 pull type bus
  dp1_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp1 glitch filter debounce clock select bus
  dp1_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp1 glitch filter bypass bus
  dp1_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp1 PES enable bus
  dp1_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp1 PES input enable bus
  dp1_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp1 PES safe value bus
  dp1_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp1 LVDS enable control bus
  dp1_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp1 input termination enable bus
  dp1_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp2 async input from pad bus
  dp2_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp2 gpio out to buf bus
  dp2_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp2 gpio out enable bus
  dp2_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp2 pinmux data to gpio bus
  dp2_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp2 pinmux enable to gpio bus
  dp2_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp2 GP DATA IN out bus
  dp2_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp2 data out to pinmux bus
  dp2_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp2 pinmux muxsel out bus
  dp2_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp2 in function enable out bus
  dp2_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp2 analog mode select bus
  dp2_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp2 drive strength 0 bus
  dp2_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp2 drive strength 1 bus
  dp2_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp2 slew control bus
  dp2_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp2 schmitt trigger bus
  dp2_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp2 mode 0 bus
  dp2_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp2 mode 1 bus
  dp2_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp2 input enable bus
  dp2_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp2 direction bus
  dp2_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp2 pull enable bus
  dp2_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp2 pull type bus
  dp2_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp2 glitch filter debounce clock select bus
  dp2_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp2 glitch filter bypass bus
  dp2_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp2 PES enable bus
  dp2_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp2 PES input enable bus
  dp2_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp2 PES safe value bus
  dp2_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp2 LVDS enable control bus
  dp2_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp2 input termination enable bus
  dp2_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp3 async input from pad bus
  dp3_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp3 gpio out to buf bus
  dp3_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp3 gpio out enable bus
  dp3_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp3 pinmux data to gpio bus
  dp3_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp3 pinmux enable to gpio bus
  dp3_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp3 GP DATA IN out bus
  dp3_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp3 data out to pinmux bus
  dp3_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp3 pinmux muxsel out bus
  dp3_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp3 in function enable out bus
  dp3_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp3 analog mode select bus
  dp3_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp3 drive strength 0 bus
  dp3_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp3 drive strength 1 bus
  dp3_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp3 slew control bus
  dp3_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp3 schmitt trigger bus
  dp3_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp3 mode 0 bus
  dp3_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp3 mode 1 bus
  dp3_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp3 input enable bus
  dp3_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp3 direction bus
  dp3_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp3 pull enable bus
  dp3_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp3 pull type bus
  dp3_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp3 glitch filter debounce clock select bus
  dp3_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp3 glitch filter bypass bus
  dp3_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp3 PES enable bus
  dp3_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp3 PES input enable bus
  dp3_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp3 PES safe value bus
  dp3_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp3 LVDS enable control bus
  dp3_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp3 input termination enable bus
  dp3_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp4 async input from pad bus
  dp4_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp4 gpio out to buf bus
  dp4_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp4 gpio out enable bus
  dp4_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp4 pinmux data to gpio bus
  dp4_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp4 pinmux enable to gpio bus
  dp4_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp4 GP DATA IN out bus
  dp4_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp4 data out to pinmux bus
  dp4_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp4 pinmux muxsel out bus
  dp4_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp4 in function enable out bus
  dp4_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp4 analog mode select bus
  dp4_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp4 drive strength 0 bus
  dp4_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp4 drive strength 1 bus
  dp4_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp4 slew control bus
  dp4_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp4 schmitt trigger bus
  dp4_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp4 mode 0 bus
  dp4_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp4 mode 1 bus
  dp4_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp4 input enable bus
  dp4_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp4 direction bus
  dp4_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp4 pull enable bus
  dp4_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp4 pull type bus
  dp4_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp4 glitch filter debounce clock select bus
  dp4_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp4 glitch filter bypass bus
  dp4_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp4 PES enable bus
  dp4_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp4 PES input enable bus
  dp4_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp4 PES safe value bus
  dp4_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp4 LVDS enable control bus
  dp4_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp4 input termination enable bus
  dp4_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp5 async input from pad bus
  dp5_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp5 gpio out to buf bus
  dp5_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp5 gpio out enable bus
  dp5_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp5 pinmux data to gpio bus
  dp5_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp5 pinmux enable to gpio bus
  dp5_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp5 GP DATA IN out bus
  dp5_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp5 data out to pinmux bus
  dp5_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp5 pinmux muxsel out bus
  dp5_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp5 in function enable out bus
  dp5_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp5 analog mode select bus
  dp5_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp5 drive strength 0 bus
  dp5_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp5 drive strength 1 bus
  dp5_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp5 slew control bus
  dp5_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp5 schmitt trigger bus
  dp5_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp5 mode 0 bus
  dp5_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp5 mode 1 bus
  dp5_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp5 input enable bus
  dp5_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp5 direction bus
  dp5_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp5 pull enable bus
  dp5_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp5 pull type bus
  dp5_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp5 glitch filter debounce clock select bus
  dp5_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp5 glitch filter bypass bus
  dp5_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp5 PES enable bus
  dp5_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp5 PES input enable bus
  dp5_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp5 PES safe value bus
  dp5_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp5 LVDS enable control bus
  dp5_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp5 input termination enable bus
  dp5_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp6 async input from pad bus
  dp6_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp6 gpio out to buf bus
  dp6_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp6 gpio out enable bus
  dp6_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp6 pinmux data to gpio bus
  dp6_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp6 pinmux enable to gpio bus
  dp6_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp6 GP DATA IN out bus
  dp6_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp6 data out to pinmux bus
  dp6_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp6 pinmux muxsel out bus
  dp6_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp6 in function enable out bus
  dp6_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp6 analog mode select bus
  dp6_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp6 drive strength 0 bus
  dp6_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp6 drive strength 1 bus
  dp6_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp6 slew control bus
  dp6_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp6 schmitt trigger bus
  dp6_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp6 mode 0 bus
  dp6_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp6 mode 1 bus
  dp6_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp6 input enable bus
  dp6_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp6 direction bus
  dp6_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp6 pull enable bus
  dp6_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp6 pull type bus
  dp6_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp6 glitch filter debounce clock select bus
  dp6_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp6 glitch filter bypass bus
  dp6_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp6 PES enable bus
  dp6_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp6 PES input enable bus
  dp6_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp6 PES safe value bus
  dp6_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp6 LVDS enable control bus
  dp6_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp6 input termination enable bus
  dp6_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // dp7 async input from pad bus
  dp7_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // dp7 gpio out to buf bus
  dp7_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // dp7 gpio out enable bus
  dp7_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // dp7 pinmux data to gpio bus
  dp7_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // dp7 pinmux enable to gpio bus
  dp7_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // dp7 GP DATA IN out bus
  dp7_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // dp7 data out to pinmux bus
  dp7_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // dp7 pinmux muxsel out bus
  dp7_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // dp7 in function enable out bus
  dp7_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // dp7 analog mode select bus
  dp7_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // dp7 drive strength 0 bus
  dp7_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // dp7 drive strength 1 bus
  dp7_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // dp7 slew control bus
  dp7_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // dp7 schmitt trigger bus
  dp7_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // dp7 mode 0 bus
  dp7_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // dp7 mode 1 bus
  dp7_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // dp7 input enable bus
  dp7_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // dp7 direction bus
  dp7_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // dp7 pull enable bus
  dp7_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // dp7 pull type bus
  dp7_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // dp7 glitch filter debounce clock select bus
  dp7_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // dp7 glitch filter bypass bus
  dp7_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // dp7 PES enable bus
  dp7_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // dp7 PES input enable bus
  dp7_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // dp7 PES safe value bus
  dp7_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // dp7 LVDS enable control bus
  dp7_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // dp7 input termination enable bus
  dp7_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // mp0 async input from pad bus
  mp0_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // mp0 gpio out to buf bus
  mp0_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // mp0 gpio out enable bus
  mp0_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // mp0 pinmux data to gpio bus
  mp0_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // mp0 pinmux enable to gpio bus
  mp0_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // mp0 GP DATA IN out bus
  mp0_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // mp0 data out to pinmux bus
  mp0_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // mp0 pinmux muxsel out bus
  mp0_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // mp0 in function enable out bus
  mp0_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // mp0 analog mode select bus
  mp0_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // mp0 drive strength 0 bus
  mp0_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // mp0 drive strength 1 bus
  mp0_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // mp0 slew control bus
  mp0_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // mp0 schmitt trigger bus
  mp0_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // mp0 mode 0 bus
  mp0_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // mp0 mode 1 bus
  mp0_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // mp0 input enable bus
  mp0_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // mp0 direction bus
  mp0_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // mp0 pull enable bus
  mp0_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // mp0 pull type bus
  mp0_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // mp0 glitch filter debounce clock select bus
  mp0_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // mp0 glitch filter bypass bus
  mp0_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // mp0 PES enable bus
  mp0_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // mp0 PES input enable bus
  mp0_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // mp0 PES safe value bus
  mp0_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // mp0 LVDS enable control bus
  mp0_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // mp0 input termination enable bus
  mp0_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // mp1 async input from pad bus
  mp1_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // mp1 gpio out to buf bus
  mp1_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // mp1 gpio out enable bus
  mp1_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // mp1 pinmux data to gpio bus
  mp1_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // mp1 pinmux enable to gpio bus
  mp1_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // mp1 GP DATA IN out bus
  mp1_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // mp1 data out to pinmux bus
  mp1_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // mp1 pinmux muxsel out bus
  mp1_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // mp1 in function enable out bus
  mp1_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // mp1 analog mode select bus
  mp1_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // mp1 drive strength 0 bus
  mp1_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // mp1 drive strength 1 bus
  mp1_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // mp1 slew control bus
  mp1_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // mp1 schmitt trigger bus
  mp1_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // mp1 mode 0 bus
  mp1_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // mp1 mode 1 bus
  mp1_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // mp1 input enable bus
  mp1_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // mp1 direction bus
  mp1_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // mp1 pull enable bus
  mp1_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // mp1 pull type bus
  mp1_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // mp1 glitch filter debounce clock select bus
  mp1_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // mp1 glitch filter bypass bus
  mp1_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // mp1 PES enable bus
  mp1_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // mp1 PES input enable bus
  mp1_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // mp1 PES safe value bus
  mp1_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // mp1 LVDS enable control bus
  mp1_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // mp1 input termination enable bus
  mp1_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // mp2 async input from pad bus
  mp2_async_in_from_pad_mscbus,                  // Bus Miscellanous Busdef

  // mp2 gpio out to buf bus
  mp2_gpio_out_2_buf_mscbus,                     // Bus Miscellanous Busdef

  // mp2 gpio out enable bus
  mp2_gpio_out_en_2_buf_mscbus,                  // Bus Miscellanous Busdef

  // mp2 pinmux data to gpio bus
  mp2_pinmuxdata_2_gpio_mscbus,                  // Bus Miscellanous Busdef

  // mp2 pinmux enable to gpio bus
  mp2_pinmuxen_2_gpio_mscbus,                    // Bus Miscellanous Busdef

  // mp2 GP DATA IN out bus
  mp2_GP_DATA_IN_out_mscbus,                     // Bus Miscellanous Busdef

  // mp2 data out to pinmux bus
  mp2_data_out_2_pinmux_mscbus,                  // Bus Miscellanous Busdef

  // mp2 pinmux muxsel out bus
  mp2_pinmux_muxsel_out_mscbus,                  // Bus Miscellanous Busdef

  // mp2 in function enable out bus
  mp2_in_function_en_out_mscbus,                 // Bus Miscellanous Busdef

  // mp2 analog mode select bus
  mp2_amsel_out_mscbus,                          // Bus Miscellanous Busdef

  // mp2 drive strength 0 bus
  mp2_ds0_out_mscbus,                            // Bus Miscellanous Busdef

  // mp2 drive strength 1 bus
  mp2_ds1_out_mscbus,                            // Bus Miscellanous Busdef

  // mp2 slew control bus
  mp2_slew_out_mscbus,                           // Bus Miscellanous Busdef

  // mp2 schmitt trigger bus
  mp2_schmitt_out_mscbus,                        // Bus Miscellanous Busdef

  // mp2 mode 0 bus
  mp2_mode0_out_mscbus,                          // Bus Miscellanous Busdef

  // mp2 mode 1 bus
  mp2_mode1_out_mscbus,                          // Bus Miscellanous Busdef

  // mp2 input enable bus
  mp2_inena_out_mscbus,                          // Bus Miscellanous Busdef

  // mp2 direction bus
  mp2_dir_out_mscbus,                            // Bus Miscellanous Busdef

  // mp2 pull enable bus
  mp2_pull_en_out_mscbus,                        // Bus Miscellanous Busdef

  // mp2 pull type bus
  mp2_pull_type_out_mscbus,                      // Bus Miscellanous Busdef

  // mp2 glitch filter debounce clock select bus
  mp2_glitch_filter_debounce_clk_sel_out_mscbus, // Bus Miscellanous Busdef

  // mp2 glitch filter bypass bus
  mp2_glitch_filter_bypass_out_mscbus,           // Bus Miscellanous Busdef

  // mp2 PES enable bus
  mp2_pes_en_out_mscbus,                         // Bus Miscellanous Busdef

  // mp2 PES input enable bus
  mp2_pes_in_en_out_mscbus,                      // Bus Miscellanous Busdef

  // mp2 PES safe value bus
  mp2_pes_safeval_out_mscbus,                    // Bus Miscellanous Busdef

  // mp2 LVDS enable control bus
  mp2_lvds_en_ctrl_out_mscbus,                   // Bus Miscellanous Busdef

  // mp2 input termination enable bus
  mp2_in_termination_en_out_mscbus,              // Bus Miscellanous Busdef

  // ap async input from pad bus
  ap_async_in_from_pad_mscbus,                   // Bus Miscellanous Busdef

  // ap gpio out to buf bus
  ap_gpio_out_2_buf_mscbus,                      // Bus Miscellanous Busdef

  // ap gpio out enable bus
  ap_gpio_out_en_2_buf_mscbus,                   // Bus Miscellanous Busdef

  // ap pinmux data to gpio bus
  ap_pinmuxdata_2_gpio_mscbus,                   // Bus Miscellanous Busdef

  // ap pinmux enable to gpio bus
  ap_pinmuxen_2_gpio_mscbus,                     // Bus Miscellanous Busdef

  // ap GP DATA IN out bus
  ap_GP_DATA_IN_out_mscbus,                      // Bus Miscellanous Busdef

  // ap data out to pinmux bus
  ap_data_out_2_pinmux_mscbus,                   // Bus Miscellanous Busdef

  // ap pinmux muxsel out bus
  ap_pinmux_muxsel_out_mscbus,                   // Bus Miscellanous Busdef

  // ap in function enable out bus
  ap_in_function_en_out_mscbus,                  // Bus Miscellanous Busdef

  // ap analog mode select bus
  ap_amsel_out_mscbus,                           // Bus Miscellanous Busdef

  // ap drive strength 0 bus
  ap_ds0_out_mscbus,                             // Bus Miscellanous Busdef

  // ap drive strength 1 bus
  ap_ds1_out_mscbus,                             // Bus Miscellanous Busdef

  // ap slew control bus
  ap_slew_out_mscbus,                            // Bus Miscellanous Busdef

  // ap schmitt trigger bus
  ap_schmitt_out_mscbus,                         // Bus Miscellanous Busdef

  // ap mode 0 bus
  ap_mode0_out_mscbus,                           // Bus Miscellanous Busdef

  // ap mode 1 bus
  ap_mode1_out_mscbus,                           // Bus Miscellanous Busdef

  // ap input enable bus
  ap_inena_out_mscbus,                           // Bus Miscellanous Busdef

  // ap direction bus
  ap_dir_out_mscbus,                             // Bus Miscellanous Busdef

  // ap pull enable bus
  ap_pull_en_out_mscbus,                         // Bus Miscellanous Busdef

  // ap pull type bus
  ap_pull_type_out_mscbus,                       // Bus Miscellanous Busdef

  // ap glitch filter debounce clock select bus
  ap_glitch_filter_debounce_clk_sel_out_mscbus,  // Bus Miscellanous Busdef

  // ap glitch filter bypass bus
  ap_glitch_filter_bypass_out_mscbus,            // Bus Miscellanous Busdef

  // ap PES enable bus
  ap_pes_en_out_mscbus,                          // Bus Miscellanous Busdef

  // ap PES input enable bus
  ap_pes_in_en_out_mscbus,                       // Bus Miscellanous Busdef

  // ap PES safe value bus
  ap_pes_safeval_out_mscbus,                     // Bus Miscellanous Busdef

  // ap LVDS enable control bus
  ap_lvds_en_ctrl_out_mscbus,                    // Bus Miscellanous Busdef

  // ap input termination enable bus
  ap_in_termination_en_out_mscbus,               // Bus Miscellanous Busdef

  // DP0_0 input mux peripheral bus
  DP0_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_1 input mux peripheral bus
  DP0_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_1 output demux peripheral bus
  DP0_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_2 input mux peripheral bus
  DP0_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_3 input mux peripheral bus
  DP0_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_3 output demux peripheral bus
  DP0_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_4 input mux peripheral bus
  DP0_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_5 input mux peripheral bus
  DP0_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_5 output demux peripheral bus
  DP0_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_6 input mux peripheral bus
  DP0_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_7 input mux peripheral bus
  DP0_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_7 output demux peripheral bus
  DP0_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_8 input mux peripheral bus
  DP0_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_8 output demux peripheral bus
  DP0_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_9 input mux peripheral bus
  DP0_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP0_9 output demux peripheral bus
  DP0_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP0_10 input mux peripheral bus
  DP0_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_11 input mux peripheral bus
  DP0_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_12 input mux peripheral bus
  DP0_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_13 input mux peripheral bus
  DP0_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_13 output demux peripheral bus
  DP0_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_14 input mux peripheral bus
  DP0_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_14 output demux peripheral bus
  DP0_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_15 input mux peripheral bus
  DP0_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_15 output demux peripheral bus
  DP0_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_16 input mux peripheral bus
  DP0_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_16 output demux peripheral bus
  DP0_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_17 input mux peripheral bus
  DP0_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_17 output demux peripheral bus
  DP0_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_18 input mux peripheral bus
  DP0_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_18 output demux peripheral bus
  DP0_18_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_19 input mux peripheral bus
  DP0_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_20 input mux peripheral bus
  DP0_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_21 input mux peripheral bus
  DP0_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_21 output demux peripheral bus
  DP0_21_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_22 input mux peripheral bus
  DP0_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_22 output demux peripheral bus
  DP0_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_23 input mux peripheral bus
  DP0_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_23 output demux peripheral bus
  DP0_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_24 input mux peripheral bus
  DP0_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_24 output demux peripheral bus
  DP0_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_25 input mux peripheral bus
  DP0_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_25 output demux peripheral bus
  DP0_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_26 input mux peripheral bus
  DP0_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_26 output demux peripheral bus
  DP0_26_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_27 input mux peripheral bus
  DP0_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_27 output demux peripheral bus
  DP0_27_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_28 input mux peripheral bus
  DP0_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_28 output demux peripheral bus
  DP0_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_29 input mux peripheral bus
  DP0_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_29 output demux peripheral bus
  DP0_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_30 input mux peripheral bus
  DP0_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_30 output demux peripheral bus
  DP0_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP0_31 input mux peripheral bus
  DP0_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP0_31 output demux peripheral bus
  DP0_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_0 input mux peripheral bus
  DP1_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_0 output demux peripheral bus
  DP1_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_1 input mux peripheral bus
  DP1_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_1 output demux peripheral bus
  DP1_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_2 input mux peripheral bus
  DP1_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_2 output demux peripheral bus
  DP1_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_3 input mux peripheral bus
  DP1_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_3 output demux peripheral bus
  DP1_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_4 input mux peripheral bus
  DP1_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_4 output demux peripheral bus
  DP1_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_5 input mux peripheral bus
  DP1_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_5 output demux peripheral bus
  DP1_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_6 input mux peripheral bus
  DP1_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_6 output demux peripheral bus
  DP1_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_7 input mux peripheral bus
  DP1_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_7 output demux peripheral bus
  DP1_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_8 input mux peripheral bus
  DP1_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_8 output demux peripheral bus
  DP1_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_9 input mux peripheral bus
  DP1_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP1_9 output demux peripheral bus
  DP1_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP1_10 input mux peripheral bus
  DP1_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_10 output demux peripheral bus
  DP1_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_11 input mux peripheral bus
  DP1_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_11 output demux peripheral bus
  DP1_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_12 input mux peripheral bus
  DP1_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_12 output demux peripheral bus
  DP1_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_13 input mux peripheral bus
  DP1_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_13 output demux peripheral bus
  DP1_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_14 input mux peripheral bus
  DP1_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_14 output demux peripheral bus
  DP1_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_15 input mux peripheral bus
  DP1_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_15 output demux peripheral bus
  DP1_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_16 input mux peripheral bus
  DP1_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_16 output demux peripheral bus
  DP1_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_17 input mux peripheral bus
  DP1_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_17 output demux peripheral bus
  DP1_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_18 input mux peripheral bus
  DP1_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_18 output demux peripheral bus
  DP1_18_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_19 input mux peripheral bus
  DP1_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_19 output demux peripheral bus
  DP1_19_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_20 input mux peripheral bus
  DP1_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_20 output demux peripheral bus
  DP1_20_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_21 input mux peripheral bus
  DP1_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_21 output demux peripheral bus
  DP1_21_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_22 input mux peripheral bus
  DP1_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_22 output demux peripheral bus
  DP1_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_23 input mux peripheral bus
  DP1_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_23 output demux peripheral bus
  DP1_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_24 input mux peripheral bus
  DP1_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_24 output demux peripheral bus
  DP1_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_25 input mux peripheral bus
  DP1_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_26 input mux peripheral bus
  DP1_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_27 input mux peripheral bus
  DP1_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_28 input mux peripheral bus
  DP1_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_28 output demux peripheral bus
  DP1_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_29 input mux peripheral bus
  DP1_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_29 output demux peripheral bus
  DP1_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_30 input mux peripheral bus
  DP1_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_30 output demux peripheral bus
  DP1_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP1_31 input mux peripheral bus
  DP1_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP1_31 output demux peripheral bus
  DP1_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_0 input mux peripheral bus
  DP2_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_0 output demux peripheral bus
  DP2_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP2_1 input mux peripheral bus
  DP2_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_2 input mux peripheral bus
  DP2_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_2 output demux peripheral bus
  DP2_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP2_3 input mux peripheral bus
  DP2_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_3 output demux peripheral bus
  DP2_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP2_4 input mux peripheral bus
  DP2_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_5 input mux peripheral bus
  DP2_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_6 input mux peripheral bus
  DP2_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_6 output demux peripheral bus
  DP2_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP2_7 input mux peripheral bus
  DP2_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_8 input mux peripheral bus
  DP2_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_9 input mux peripheral bus
  DP2_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP2_10 input mux peripheral bus
  DP2_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_11 input mux peripheral bus
  DP2_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_12 input mux peripheral bus
  DP2_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_12 output demux peripheral bus
  DP2_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_13 input mux peripheral bus
  DP2_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_13 output demux peripheral bus
  DP2_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_14 input mux peripheral bus
  DP2_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_15 input mux peripheral bus
  DP2_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_15 output demux peripheral bus
  DP2_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_16 input mux peripheral bus
  DP2_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_16 output demux peripheral bus
  DP2_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_17 input mux peripheral bus
  DP2_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_17 output demux peripheral bus
  DP2_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_18 input mux peripheral bus
  DP2_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_19 input mux peripheral bus
  DP2_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_20 input mux peripheral bus
  DP2_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_20 output demux peripheral bus
  DP2_20_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_21 input mux peripheral bus
  DP2_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_22 input mux peripheral bus
  DP2_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_22 output demux peripheral bus
  DP2_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_23 input mux peripheral bus
  DP2_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_23 output demux peripheral bus
  DP2_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_24 input mux peripheral bus
  DP2_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_24 output demux peripheral bus
  DP2_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_25 input mux peripheral bus
  DP2_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_26 input mux peripheral bus
  DP2_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_26 output demux peripheral bus
  DP2_26_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_27 input mux peripheral bus
  DP2_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_27 output demux peripheral bus
  DP2_27_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_28 input mux peripheral bus
  DP2_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_28 output demux peripheral bus
  DP2_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_29 input mux peripheral bus
  DP2_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_29 output demux peripheral bus
  DP2_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_30 input mux peripheral bus
  DP2_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_30 output demux peripheral bus
  DP2_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP2_31 input mux peripheral bus
  DP2_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP2_31 output demux peripheral bus
  DP2_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_0 input mux peripheral bus
  DP3_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_0 output demux peripheral bus
  DP3_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_1 input mux peripheral bus
  DP3_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_1 output demux peripheral bus
  DP3_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_2 input mux peripheral bus
  DP3_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_2 output demux peripheral bus
  DP3_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_3 input mux peripheral bus
  DP3_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_3 output demux peripheral bus
  DP3_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_4 input mux peripheral bus
  DP3_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_4 output demux peripheral bus
  DP3_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_5 input mux peripheral bus
  DP3_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_5 output demux peripheral bus
  DP3_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_6 input mux peripheral bus
  DP3_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_6 output demux peripheral bus
  DP3_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_7 input mux peripheral bus
  DP3_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_7 output demux peripheral bus
  DP3_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_8 input mux peripheral bus
  DP3_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_8 output demux peripheral bus
  DP3_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_9 input mux peripheral bus
  DP3_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP3_9 output demux peripheral bus
  DP3_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP3_10 input mux peripheral bus
  DP3_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_10 output demux peripheral bus
  DP3_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_11 input mux peripheral bus
  DP3_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_11 output demux peripheral bus
  DP3_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_12 input mux peripheral bus
  DP3_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_13 input mux peripheral bus
  DP3_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_13 output demux peripheral bus
  DP3_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_14 input mux peripheral bus
  DP3_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_15 input mux peripheral bus
  DP3_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_15 output demux peripheral bus
  DP3_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_16 input mux peripheral bus
  DP3_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_16 output demux peripheral bus
  DP3_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_17 input mux peripheral bus
  DP3_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_17 output demux peripheral bus
  DP3_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_18 input mux peripheral bus
  DP3_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_19 input mux peripheral bus
  DP3_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_20 input mux peripheral bus
  DP3_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_21 input mux peripheral bus
  DP3_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_22 input mux peripheral bus
  DP3_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_23 input mux peripheral bus
  DP3_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_24 input mux peripheral bus
  DP3_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_24 output demux peripheral bus
  DP3_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_25 input mux peripheral bus
  DP3_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_25 output demux peripheral bus
  DP3_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_26 input mux peripheral bus
  DP3_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_26 output demux peripheral bus
  DP3_26_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_27 input mux peripheral bus
  DP3_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_27 output demux peripheral bus
  DP3_27_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_28 input mux peripheral bus
  DP3_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_28 output demux peripheral bus
  DP3_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_29 input mux peripheral bus
  DP3_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_30 input mux peripheral bus
  DP3_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_30 output demux peripheral bus
  DP3_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP3_31 input mux peripheral bus
  DP3_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP3_31 output demux peripheral bus
  DP3_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_0 input mux peripheral bus
  DP4_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_0 output demux peripheral bus
  DP4_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_1 input mux peripheral bus
  DP4_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_1 output demux peripheral bus
  DP4_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_2 input mux peripheral bus
  DP4_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_2 output demux peripheral bus
  DP4_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_3 input mux peripheral bus
  DP4_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_3 output demux peripheral bus
  DP4_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_4 input mux peripheral bus
  DP4_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_4 output demux peripheral bus
  DP4_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_5 input mux peripheral bus
  DP4_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_6 input mux peripheral bus
  DP4_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_6 output demux peripheral bus
  DP4_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_7 input mux peripheral bus
  DP4_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_7 output demux peripheral bus
  DP4_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_8 input mux peripheral bus
  DP4_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_9 input mux peripheral bus
  DP4_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP4_9 output demux peripheral bus
  DP4_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP4_10 input mux peripheral bus
  DP4_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_10 output demux peripheral bus
  DP4_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_11 input mux peripheral bus
  DP4_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_11 output demux peripheral bus
  DP4_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_12 input mux peripheral bus
  DP4_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_12 output demux peripheral bus
  DP4_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_13 input mux peripheral bus
  DP4_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_13 output demux peripheral bus
  DP4_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_14 input mux peripheral bus
  DP4_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_14 output demux peripheral bus
  DP4_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_15 input mux peripheral bus
  DP4_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_15 output demux peripheral bus
  DP4_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_16 input mux peripheral bus
  DP4_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_16 output demux peripheral bus
  DP4_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_17 input mux peripheral bus
  DP4_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_17 output demux peripheral bus
  DP4_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_18 input mux peripheral bus
  DP4_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_18 output demux peripheral bus
  DP4_18_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_19 input mux peripheral bus
  DP4_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_20 input mux peripheral bus
  DP4_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_21 input mux peripheral bus
  DP4_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_22 input mux peripheral bus
  DP4_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_22 output demux peripheral bus
  DP4_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_23 input mux peripheral bus
  DP4_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_24 input mux peripheral bus
  DP4_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_25 input mux peripheral bus
  DP4_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_25 output demux peripheral bus
  DP4_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_26 input mux peripheral bus
  DP4_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_27 input mux peripheral bus
  DP4_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_27 output demux peripheral bus
  DP4_27_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_28 input mux peripheral bus
  DP4_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_28 output demux peripheral bus
  DP4_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_29 input mux peripheral bus
  DP4_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_29 output demux peripheral bus
  DP4_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_30 input mux peripheral bus
  DP4_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_30 output demux peripheral bus
  DP4_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP4_31 input mux peripheral bus
  DP4_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP4_31 output demux peripheral bus
  DP4_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_0 input mux peripheral bus
  DP5_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_1 input mux peripheral bus
  DP5_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_1 output demux peripheral bus
  DP5_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_2 input mux peripheral bus
  DP5_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_2 output demux peripheral bus
  DP5_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_3 input mux peripheral bus
  DP5_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_3 output demux peripheral bus
  DP5_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_4 input mux peripheral bus
  DP5_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_4 output demux peripheral bus
  DP5_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_5 input mux peripheral bus
  DP5_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_5 output demux peripheral bus
  DP5_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_6 input mux peripheral bus
  DP5_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_6 output demux peripheral bus
  DP5_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_7 input mux peripheral bus
  DP5_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_8 input mux peripheral bus
  DP5_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_8 output demux peripheral bus
  DP5_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_9 input mux peripheral bus
  DP5_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP5_9 output demux peripheral bus
  DP5_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP5_10 input mux peripheral bus
  DP5_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_10 output demux peripheral bus
  DP5_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_11 input mux peripheral bus
  DP5_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_11 output demux peripheral bus
  DP5_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_12 input mux peripheral bus
  DP5_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_12 output demux peripheral bus
  DP5_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_13 input mux peripheral bus
  DP5_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_13 output demux peripheral bus
  DP5_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_14 input mux peripheral bus
  DP5_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_15 input mux peripheral bus
  DP5_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_15 output demux peripheral bus
  DP5_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_16 input mux peripheral bus
  DP5_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_16 output demux peripheral bus
  DP5_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_17 input mux peripheral bus
  DP5_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_17 output demux peripheral bus
  DP5_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_18 input mux peripheral bus
  DP5_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_19 input mux peripheral bus
  DP5_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_19 output demux peripheral bus
  DP5_19_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_20 input mux peripheral bus
  DP5_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_21 input mux peripheral bus
  DP5_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_21 output demux peripheral bus
  DP5_21_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_22 input mux peripheral bus
  DP5_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_22 output demux peripheral bus
  DP5_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_23 input mux peripheral bus
  DP5_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_23 output demux peripheral bus
  DP5_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_24 input mux peripheral bus
  DP5_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_24 output demux peripheral bus
  DP5_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_25 input mux peripheral bus
  DP5_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_25 output demux peripheral bus
  DP5_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_26 input mux peripheral bus
  DP5_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_26 output demux peripheral bus
  DP5_26_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_27 input mux peripheral bus
  DP5_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_28 input mux peripheral bus
  DP5_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_28 output demux peripheral bus
  DP5_28_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_29 input mux peripheral bus
  DP5_29_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_29 output demux peripheral bus
  DP5_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_30 input mux peripheral bus
  DP5_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_30 output demux peripheral bus
  DP5_30_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP5_31 input mux peripheral bus
  DP5_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP5_31 output demux peripheral bus
  DP5_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_0 input mux peripheral bus
  DP6_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_0 output demux peripheral bus
  DP6_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_1 input mux peripheral bus
  DP6_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_1 output demux peripheral bus
  DP6_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_2 input mux peripheral bus
  DP6_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_2 output demux peripheral bus
  DP6_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_3 input mux peripheral bus
  DP6_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_3 output demux peripheral bus
  DP6_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_4 input mux peripheral bus
  DP6_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_4 output demux peripheral bus
  DP6_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_5 input mux peripheral bus
  DP6_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_5 output demux peripheral bus
  DP6_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_6 input mux peripheral bus
  DP6_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_6 output demux peripheral bus
  DP6_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_7 input mux peripheral bus
  DP6_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_7 output demux peripheral bus
  DP6_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_8 input mux peripheral bus
  DP6_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_8 output demux peripheral bus
  DP6_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_9 input mux peripheral bus
  DP6_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP6_9 output demux peripheral bus
  DP6_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP6_10 input mux peripheral bus
  DP6_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_10 output demux peripheral bus
  DP6_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_11 input mux peripheral bus
  DP6_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_12 input mux peripheral bus
  DP6_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_12 output demux peripheral bus
  DP6_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_13 input mux peripheral bus
  DP6_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_13 output demux peripheral bus
  DP6_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_14 input mux peripheral bus
  DP6_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_14 output demux peripheral bus
  DP6_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_15 input mux peripheral bus
  DP6_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_15 output demux peripheral bus
  DP6_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_16 input mux peripheral bus
  DP6_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_16 output demux peripheral bus
  DP6_16_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_17 input mux peripheral bus
  DP6_17_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_18 input mux peripheral bus
  DP6_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_18 output demux peripheral bus
  DP6_18_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_19 input mux peripheral bus
  DP6_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_19 output demux peripheral bus
  DP6_19_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_20 input mux peripheral bus
  DP6_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_21 input mux peripheral bus
  DP6_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_21 output demux peripheral bus
  DP6_21_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_22 input mux peripheral bus
  DP6_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_22 output demux peripheral bus
  DP6_22_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_23 input mux peripheral bus
  DP6_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_23 output demux peripheral bus
  DP6_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_24 input mux peripheral bus
  DP6_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_24 output demux peripheral bus
  DP6_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_25 input mux peripheral bus
  DP6_25_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_25 output demux peripheral bus
  DP6_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP6_26 input mux peripheral bus
  DP6_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP6_27 input mux peripheral bus
  DP6_27_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_0 input mux peripheral bus
  DP7_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_1 input mux peripheral bus
  DP7_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_1 output demux peripheral bus
  DP7_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP7_2 input mux peripheral bus
  DP7_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_3 input mux peripheral bus
  DP7_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_4 input mux peripheral bus
  DP7_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_5 input mux peripheral bus
  DP7_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_6 input mux peripheral bus
  DP7_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_6 output demux peripheral bus
  DP7_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP7_7 input mux peripheral bus
  DP7_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_7 output demux peripheral bus
  DP7_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP7_8 input mux peripheral bus
  DP7_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_8 output demux peripheral bus
  DP7_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP7_9 input mux peripheral bus
  DP7_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // DP7_9 output demux peripheral bus
  DP7_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // DP7_10 input mux peripheral bus
  DP7_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_10 output demux peripheral bus
  DP7_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP7_11 input mux peripheral bus
  DP7_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_11 output demux peripheral bus
  DP7_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP7_12 input mux peripheral bus
  DP7_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_12 output demux peripheral bus
  DP7_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP7_13 input mux peripheral bus
  DP7_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_13 output demux peripheral bus
  DP7_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP7_14 input mux peripheral bus
  DP7_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_14 output demux peripheral bus
  DP7_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // DP7_15 input mux peripheral bus
  DP7_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // DP7_15 output demux peripheral bus
  DP7_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_0 input mux peripheral bus
  MP0_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_0 output demux peripheral bus
  MP0_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_1 input mux peripheral bus
  MP0_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_1 output demux peripheral bus
  MP0_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_2 input mux peripheral bus
  MP0_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_2 output demux peripheral bus
  MP0_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_3 input mux peripheral bus
  MP0_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_3 output demux peripheral bus
  MP0_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_4 input mux peripheral bus
  MP0_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_4 output demux peripheral bus
  MP0_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_5 output demux peripheral bus
  MP0_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_6 input mux peripheral bus
  MP0_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_6 output demux peripheral bus
  MP0_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_7 input mux peripheral bus
  MP0_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_7 output demux peripheral bus
  MP0_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_8 input mux peripheral bus
  MP0_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_8 output demux peripheral bus
  MP0_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_9 input mux peripheral bus
  MP0_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP0_9 output demux peripheral bus
  MP0_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP0_10 input mux peripheral bus
  MP0_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_10 output demux peripheral bus
  MP0_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_11 output demux peripheral bus
  MP0_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_12 input mux peripheral bus
  MP0_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_12 output demux peripheral bus
  MP0_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_13 input mux peripheral bus
  MP0_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_13 output demux peripheral bus
  MP0_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_14 input mux peripheral bus
  MP0_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_15 input mux peripheral bus
  MP0_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_15 output demux peripheral bus
  MP0_15_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_16 input mux peripheral bus
  MP0_16_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_17 output demux peripheral bus
  MP0_17_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_18 input mux peripheral bus
  MP0_18_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_19 input mux peripheral bus
  MP0_19_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_19 output demux peripheral bus
  MP0_19_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_20 input mux peripheral bus
  MP0_20_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_21 input mux peripheral bus
  MP0_21_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_21 output demux peripheral bus
  MP0_21_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_22 input mux peripheral bus
  MP0_22_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_23 input mux peripheral bus
  MP0_23_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_23 output demux peripheral bus
  MP0_23_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_24 input mux peripheral bus
  MP0_24_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_24 output demux peripheral bus
  MP0_24_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_25 output demux peripheral bus
  MP0_25_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_26 input mux peripheral bus
  MP0_26_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_26 output demux peripheral bus
  MP0_26_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_27 output demux peripheral bus
  MP0_27_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_28 input mux peripheral bus
  MP0_28_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_29 output demux peripheral bus
  MP0_29_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP0_30 input mux peripheral bus
  MP0_30_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_31 input mux peripheral bus
  MP0_31_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP0_31 output demux peripheral bus
  MP0_31_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP1_0 input mux peripheral bus
  MP1_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_1 input mux peripheral bus
  MP1_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_1 output demux peripheral bus
  MP1_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_2 input mux peripheral bus
  MP1_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_2 output demux peripheral bus
  MP1_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_3 output demux peripheral bus
  MP1_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_4 input mux peripheral bus
  MP1_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_4 output demux peripheral bus
  MP1_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_5 input mux peripheral bus
  MP1_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_5 output demux peripheral bus
  MP1_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_6 input mux peripheral bus
  MP1_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_6 output demux peripheral bus
  MP1_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_7 input mux peripheral bus
  MP1_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_7 output demux peripheral bus
  MP1_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_8 input mux peripheral bus
  MP1_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_8 output demux peripheral bus
  MP1_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_9 input mux peripheral bus
  MP1_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP1_9 output demux peripheral bus
  MP1_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP1_10 input mux peripheral bus
  MP1_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP1_11 input mux peripheral bus
  MP1_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP1_12 input mux peripheral bus
  MP1_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP1_13 input mux peripheral bus
  MP1_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP1_14 input mux peripheral bus
  MP1_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP1_15 input mux peripheral bus
  MP1_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_0 input mux peripheral bus
  MP2_0_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_0 output demux peripheral bus
  MP2_0_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_1 input mux peripheral bus
  MP2_1_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_1 output demux peripheral bus
  MP2_1_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_2 input mux peripheral bus
  MP2_2_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_2 output demux peripheral bus
  MP2_2_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_3 input mux peripheral bus
  MP2_3_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_3 output demux peripheral bus
  MP2_3_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_4 input mux peripheral bus
  MP2_4_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_4 output demux peripheral bus
  MP2_4_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_5 input mux peripheral bus
  MP2_5_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_5 output demux peripheral bus
  MP2_5_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_6 input mux peripheral bus
  MP2_6_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_6 output demux peripheral bus
  MP2_6_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_7 input mux peripheral bus
  MP2_7_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_7 output demux peripheral bus
  MP2_7_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_8 input mux peripheral bus
  MP2_8_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_8 output demux peripheral bus
  MP2_8_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_9 input mux peripheral bus
  MP2_9_in_mux_peripheral_mscbus,                // Bus Miscellanous Busdef

  // MP2_9 output demux peripheral bus
  MP2_9_out_demux_peripheral_mscbus,             // Bus Miscellanous Busdef

  // MP2_10 input mux peripheral bus
  MP2_10_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_10 output demux peripheral bus
  MP2_10_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP2_11 input mux peripheral bus
  MP2_11_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_11 output demux peripheral bus
  MP2_11_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP2_12 input mux peripheral bus
  MP2_12_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_12 output demux peripheral bus
  MP2_12_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP2_13 input mux peripheral bus
  MP2_13_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_13 output demux peripheral bus
  MP2_13_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP2_14 input mux peripheral bus
  MP2_14_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_14 output demux peripheral bus
  MP2_14_out_demux_peripheral_mscbus,            // Bus Miscellanous Busdef

  // MP2_15 input mux peripheral bus
  MP2_15_in_mux_peripheral_mscbus,               // Bus Miscellanous Busdef

  // MP2_15 output demux peripheral bus
  MP2_15_out_demux_peripheral_mscbus             // Bus Miscellanous Busdef
);

// Default Interface

// dp0 async input from pad bus
output      [31:0] dp0_async_in_from_pad_mscbus;

// dp0 gpio out to buf bus
input       [31:0] dp0_gpio_out_2_buf_mscbus;

// dp0 gpio out enable bus
input       [31:0] dp0_gpio_out_en_2_buf_mscbus;

// dp0 pinmux data to gpio bus
input       [31:0] dp0_pinmuxdata_2_gpio_mscbus;

// dp0 pinmux enable to gpio bus
input       [31:0] dp0_pinmuxen_2_gpio_mscbus;

// dp0 GP DATA IN out bus
output      [31:0] dp0_GP_DATA_IN_out_mscbus;

// dp0 data out to pinmux bus
output      [31:0] dp0_data_out_2_pinmux_mscbus;

// dp0 pinmux muxsel out bus
input      [159:0] dp0_pinmux_muxsel_out_mscbus;

// dp0 in function enable out bus
input     [1023:0] dp0_in_function_en_out_mscbus;

// dp0 analog mode select bus
input       [31:0] dp0_amsel_out_mscbus;

// dp0 drive strength 0 bus
input       [31:0] dp0_ds0_out_mscbus;

// dp0 drive strength 1 bus
input       [31:0] dp0_ds1_out_mscbus;

// dp0 slew control bus
input       [31:0] dp0_slew_out_mscbus;

// dp0 schmitt trigger bus
input       [31:0] dp0_schmitt_out_mscbus;

// dp0 mode 0 bus
input       [31:0] dp0_mode0_out_mscbus;

// dp0 mode 1 bus
input       [31:0] dp0_mode1_out_mscbus;

// dp0 input enable bus
input       [31:0] dp0_inena_out_mscbus;

// dp0 direction bus
input       [31:0] dp0_dir_out_mscbus;

// dp0 pull enable bus
input       [31:0] dp0_pull_en_out_mscbus;

// dp0 pull type bus
input       [31:0] dp0_pull_type_out_mscbus;

// dp0 glitch filter debounce clock select bus
input       [63:0] dp0_glitch_filter_debounce_clk_sel_out_mscbus;

// dp0 glitch filter bypass bus
input       [31:0] dp0_glitch_filter_bypass_out_mscbus;

// dp0 PES enable bus
input      [255:0] dp0_pes_en_out_mscbus;

// dp0 PES input enable bus
input       [31:0] dp0_pes_in_en_out_mscbus;

// dp0 PES safe value bus
input       [63:0] dp0_pes_safeval_out_mscbus;

// dp0 LVDS enable control bus
input       [31:0] dp0_lvds_en_ctrl_out_mscbus;

// dp0 input termination enable bus
input       [31:0] dp0_in_termination_en_out_mscbus;

// dp1 async input from pad bus
output      [31:0] dp1_async_in_from_pad_mscbus;

// dp1 gpio out to buf bus
input       [31:0] dp1_gpio_out_2_buf_mscbus;

// dp1 gpio out enable bus
input       [31:0] dp1_gpio_out_en_2_buf_mscbus;

// dp1 pinmux data to gpio bus
input       [31:0] dp1_pinmuxdata_2_gpio_mscbus;

// dp1 pinmux enable to gpio bus
input       [31:0] dp1_pinmuxen_2_gpio_mscbus;

// dp1 GP DATA IN out bus
output      [31:0] dp1_GP_DATA_IN_out_mscbus;

// dp1 data out to pinmux bus
output      [31:0] dp1_data_out_2_pinmux_mscbus;

// dp1 pinmux muxsel out bus
input      [159:0] dp1_pinmux_muxsel_out_mscbus;

// dp1 in function enable out bus
input     [1023:0] dp1_in_function_en_out_mscbus;

// dp1 analog mode select bus
input       [31:0] dp1_amsel_out_mscbus;

// dp1 drive strength 0 bus
input       [31:0] dp1_ds0_out_mscbus;

// dp1 drive strength 1 bus
input       [31:0] dp1_ds1_out_mscbus;

// dp1 slew control bus
input       [31:0] dp1_slew_out_mscbus;

// dp1 schmitt trigger bus
input       [31:0] dp1_schmitt_out_mscbus;

// dp1 mode 0 bus
input       [31:0] dp1_mode0_out_mscbus;

// dp1 mode 1 bus
input       [31:0] dp1_mode1_out_mscbus;

// dp1 input enable bus
input       [31:0] dp1_inena_out_mscbus;

// dp1 direction bus
input       [31:0] dp1_dir_out_mscbus;

// dp1 pull enable bus
input       [31:0] dp1_pull_en_out_mscbus;

// dp1 pull type bus
input       [31:0] dp1_pull_type_out_mscbus;

// dp1 glitch filter debounce clock select bus
input       [63:0] dp1_glitch_filter_debounce_clk_sel_out_mscbus;

// dp1 glitch filter bypass bus
input       [31:0] dp1_glitch_filter_bypass_out_mscbus;

// dp1 PES enable bus
input      [255:0] dp1_pes_en_out_mscbus;

// dp1 PES input enable bus
input       [31:0] dp1_pes_in_en_out_mscbus;

// dp1 PES safe value bus
input       [63:0] dp1_pes_safeval_out_mscbus;

// dp1 LVDS enable control bus
input       [31:0] dp1_lvds_en_ctrl_out_mscbus;

// dp1 input termination enable bus
input       [31:0] dp1_in_termination_en_out_mscbus;

// dp2 async input from pad bus
output      [31:0] dp2_async_in_from_pad_mscbus;

// dp2 gpio out to buf bus
input       [31:0] dp2_gpio_out_2_buf_mscbus;

// dp2 gpio out enable bus
input       [31:0] dp2_gpio_out_en_2_buf_mscbus;

// dp2 pinmux data to gpio bus
input       [31:0] dp2_pinmuxdata_2_gpio_mscbus;

// dp2 pinmux enable to gpio bus
input       [31:0] dp2_pinmuxen_2_gpio_mscbus;

// dp2 GP DATA IN out bus
output      [31:0] dp2_GP_DATA_IN_out_mscbus;

// dp2 data out to pinmux bus
output      [31:0] dp2_data_out_2_pinmux_mscbus;

// dp2 pinmux muxsel out bus
input      [159:0] dp2_pinmux_muxsel_out_mscbus;

// dp2 in function enable out bus
input     [1023:0] dp2_in_function_en_out_mscbus;

// dp2 analog mode select bus
input       [31:0] dp2_amsel_out_mscbus;

// dp2 drive strength 0 bus
input       [31:0] dp2_ds0_out_mscbus;

// dp2 drive strength 1 bus
input       [31:0] dp2_ds1_out_mscbus;

// dp2 slew control bus
input       [31:0] dp2_slew_out_mscbus;

// dp2 schmitt trigger bus
input       [31:0] dp2_schmitt_out_mscbus;

// dp2 mode 0 bus
input       [31:0] dp2_mode0_out_mscbus;

// dp2 mode 1 bus
input       [31:0] dp2_mode1_out_mscbus;

// dp2 input enable bus
input       [31:0] dp2_inena_out_mscbus;

// dp2 direction bus
input       [31:0] dp2_dir_out_mscbus;

// dp2 pull enable bus
input       [31:0] dp2_pull_en_out_mscbus;

// dp2 pull type bus
input       [31:0] dp2_pull_type_out_mscbus;

// dp2 glitch filter debounce clock select bus
input       [63:0] dp2_glitch_filter_debounce_clk_sel_out_mscbus;

// dp2 glitch filter bypass bus
input       [31:0] dp2_glitch_filter_bypass_out_mscbus;

// dp2 PES enable bus
input      [255:0] dp2_pes_en_out_mscbus;

// dp2 PES input enable bus
input       [31:0] dp2_pes_in_en_out_mscbus;

// dp2 PES safe value bus
input       [63:0] dp2_pes_safeval_out_mscbus;

// dp2 LVDS enable control bus
input       [31:0] dp2_lvds_en_ctrl_out_mscbus;

// dp2 input termination enable bus
input       [31:0] dp2_in_termination_en_out_mscbus;

// dp3 async input from pad bus
output      [31:0] dp3_async_in_from_pad_mscbus;

// dp3 gpio out to buf bus
input       [31:0] dp3_gpio_out_2_buf_mscbus;

// dp3 gpio out enable bus
input       [31:0] dp3_gpio_out_en_2_buf_mscbus;

// dp3 pinmux data to gpio bus
input       [31:0] dp3_pinmuxdata_2_gpio_mscbus;

// dp3 pinmux enable to gpio bus
input       [31:0] dp3_pinmuxen_2_gpio_mscbus;

// dp3 GP DATA IN out bus
output      [31:0] dp3_GP_DATA_IN_out_mscbus;

// dp3 data out to pinmux bus
output      [31:0] dp3_data_out_2_pinmux_mscbus;

// dp3 pinmux muxsel out bus
input      [159:0] dp3_pinmux_muxsel_out_mscbus;

// dp3 in function enable out bus
input     [1023:0] dp3_in_function_en_out_mscbus;

// dp3 analog mode select bus
input       [31:0] dp3_amsel_out_mscbus;

// dp3 drive strength 0 bus
input       [31:0] dp3_ds0_out_mscbus;

// dp3 drive strength 1 bus
input       [31:0] dp3_ds1_out_mscbus;

// dp3 slew control bus
input       [31:0] dp3_slew_out_mscbus;

// dp3 schmitt trigger bus
input       [31:0] dp3_schmitt_out_mscbus;

// dp3 mode 0 bus
input       [31:0] dp3_mode0_out_mscbus;

// dp3 mode 1 bus
input       [31:0] dp3_mode1_out_mscbus;

// dp3 input enable bus
input       [31:0] dp3_inena_out_mscbus;

// dp3 direction bus
input       [31:0] dp3_dir_out_mscbus;

// dp3 pull enable bus
input       [31:0] dp3_pull_en_out_mscbus;

// dp3 pull type bus
input       [31:0] dp3_pull_type_out_mscbus;

// dp3 glitch filter debounce clock select bus
input       [63:0] dp3_glitch_filter_debounce_clk_sel_out_mscbus;

// dp3 glitch filter bypass bus
input       [31:0] dp3_glitch_filter_bypass_out_mscbus;

// dp3 PES enable bus
input      [255:0] dp3_pes_en_out_mscbus;

// dp3 PES input enable bus
input       [31:0] dp3_pes_in_en_out_mscbus;

// dp3 PES safe value bus
input       [63:0] dp3_pes_safeval_out_mscbus;

// dp3 LVDS enable control bus
input       [31:0] dp3_lvds_en_ctrl_out_mscbus;

// dp3 input termination enable bus
input       [31:0] dp3_in_termination_en_out_mscbus;

// dp4 async input from pad bus
output      [31:0] dp4_async_in_from_pad_mscbus;

// dp4 gpio out to buf bus
input       [31:0] dp4_gpio_out_2_buf_mscbus;

// dp4 gpio out enable bus
input       [31:0] dp4_gpio_out_en_2_buf_mscbus;

// dp4 pinmux data to gpio bus
input       [31:0] dp4_pinmuxdata_2_gpio_mscbus;

// dp4 pinmux enable to gpio bus
input       [31:0] dp4_pinmuxen_2_gpio_mscbus;

// dp4 GP DATA IN out bus
output      [31:0] dp4_GP_DATA_IN_out_mscbus;

// dp4 data out to pinmux bus
output      [31:0] dp4_data_out_2_pinmux_mscbus;

// dp4 pinmux muxsel out bus
input      [159:0] dp4_pinmux_muxsel_out_mscbus;

// dp4 in function enable out bus
input     [1023:0] dp4_in_function_en_out_mscbus;

// dp4 analog mode select bus
input       [31:0] dp4_amsel_out_mscbus;

// dp4 drive strength 0 bus
input       [31:0] dp4_ds0_out_mscbus;

// dp4 drive strength 1 bus
input       [31:0] dp4_ds1_out_mscbus;

// dp4 slew control bus
input       [31:0] dp4_slew_out_mscbus;

// dp4 schmitt trigger bus
input       [31:0] dp4_schmitt_out_mscbus;

// dp4 mode 0 bus
input       [31:0] dp4_mode0_out_mscbus;

// dp4 mode 1 bus
input       [31:0] dp4_mode1_out_mscbus;

// dp4 input enable bus
input       [31:0] dp4_inena_out_mscbus;

// dp4 direction bus
input       [31:0] dp4_dir_out_mscbus;

// dp4 pull enable bus
input       [31:0] dp4_pull_en_out_mscbus;

// dp4 pull type bus
input       [31:0] dp4_pull_type_out_mscbus;

// dp4 glitch filter debounce clock select bus
input       [63:0] dp4_glitch_filter_debounce_clk_sel_out_mscbus;

// dp4 glitch filter bypass bus
input       [31:0] dp4_glitch_filter_bypass_out_mscbus;

// dp4 PES enable bus
input      [255:0] dp4_pes_en_out_mscbus;

// dp4 PES input enable bus
input       [31:0] dp4_pes_in_en_out_mscbus;

// dp4 PES safe value bus
input       [63:0] dp4_pes_safeval_out_mscbus;

// dp4 LVDS enable control bus
input       [31:0] dp4_lvds_en_ctrl_out_mscbus;

// dp4 input termination enable bus
input       [31:0] dp4_in_termination_en_out_mscbus;

// dp5 async input from pad bus
output      [31:0] dp5_async_in_from_pad_mscbus;

// dp5 gpio out to buf bus
input       [31:0] dp5_gpio_out_2_buf_mscbus;

// dp5 gpio out enable bus
input       [31:0] dp5_gpio_out_en_2_buf_mscbus;

// dp5 pinmux data to gpio bus
input       [31:0] dp5_pinmuxdata_2_gpio_mscbus;

// dp5 pinmux enable to gpio bus
input       [31:0] dp5_pinmuxen_2_gpio_mscbus;

// dp5 GP DATA IN out bus
output      [31:0] dp5_GP_DATA_IN_out_mscbus;

// dp5 data out to pinmux bus
output      [31:0] dp5_data_out_2_pinmux_mscbus;

// dp5 pinmux muxsel out bus
input      [159:0] dp5_pinmux_muxsel_out_mscbus;

// dp5 in function enable out bus
input     [1023:0] dp5_in_function_en_out_mscbus;

// dp5 analog mode select bus
input       [31:0] dp5_amsel_out_mscbus;

// dp5 drive strength 0 bus
input       [31:0] dp5_ds0_out_mscbus;

// dp5 drive strength 1 bus
input       [31:0] dp5_ds1_out_mscbus;

// dp5 slew control bus
input       [31:0] dp5_slew_out_mscbus;

// dp5 schmitt trigger bus
input       [31:0] dp5_schmitt_out_mscbus;

// dp5 mode 0 bus
input       [31:0] dp5_mode0_out_mscbus;

// dp5 mode 1 bus
input       [31:0] dp5_mode1_out_mscbus;

// dp5 input enable bus
input       [31:0] dp5_inena_out_mscbus;

// dp5 direction bus
input       [31:0] dp5_dir_out_mscbus;

// dp5 pull enable bus
input       [31:0] dp5_pull_en_out_mscbus;

// dp5 pull type bus
input       [31:0] dp5_pull_type_out_mscbus;

// dp5 glitch filter debounce clock select bus
input       [63:0] dp5_glitch_filter_debounce_clk_sel_out_mscbus;

// dp5 glitch filter bypass bus
input       [31:0] dp5_glitch_filter_bypass_out_mscbus;

// dp5 PES enable bus
input      [255:0] dp5_pes_en_out_mscbus;

// dp5 PES input enable bus
input       [31:0] dp5_pes_in_en_out_mscbus;

// dp5 PES safe value bus
input       [63:0] dp5_pes_safeval_out_mscbus;

// dp5 LVDS enable control bus
input       [31:0] dp5_lvds_en_ctrl_out_mscbus;

// dp5 input termination enable bus
input       [31:0] dp5_in_termination_en_out_mscbus;

// dp6 async input from pad bus
output      [31:0] dp6_async_in_from_pad_mscbus;

// dp6 gpio out to buf bus
input       [31:0] dp6_gpio_out_2_buf_mscbus;

// dp6 gpio out enable bus
input       [31:0] dp6_gpio_out_en_2_buf_mscbus;

// dp6 pinmux data to gpio bus
input       [31:0] dp6_pinmuxdata_2_gpio_mscbus;

// dp6 pinmux enable to gpio bus
input       [31:0] dp6_pinmuxen_2_gpio_mscbus;

// dp6 GP DATA IN out bus
output      [31:0] dp6_GP_DATA_IN_out_mscbus;

// dp6 data out to pinmux bus
output      [31:0] dp6_data_out_2_pinmux_mscbus;

// dp6 pinmux muxsel out bus
input      [159:0] dp6_pinmux_muxsel_out_mscbus;

// dp6 in function enable out bus
input     [1023:0] dp6_in_function_en_out_mscbus;

// dp6 analog mode select bus
input       [31:0] dp6_amsel_out_mscbus;

// dp6 drive strength 0 bus
input       [31:0] dp6_ds0_out_mscbus;

// dp6 drive strength 1 bus
input       [31:0] dp6_ds1_out_mscbus;

// dp6 slew control bus
input       [31:0] dp6_slew_out_mscbus;

// dp6 schmitt trigger bus
input       [31:0] dp6_schmitt_out_mscbus;

// dp6 mode 0 bus
input       [31:0] dp6_mode0_out_mscbus;

// dp6 mode 1 bus
input       [31:0] dp6_mode1_out_mscbus;

// dp6 input enable bus
input       [31:0] dp6_inena_out_mscbus;

// dp6 direction bus
input       [31:0] dp6_dir_out_mscbus;

// dp6 pull enable bus
input       [31:0] dp6_pull_en_out_mscbus;

// dp6 pull type bus
input       [31:0] dp6_pull_type_out_mscbus;

// dp6 glitch filter debounce clock select bus
input       [63:0] dp6_glitch_filter_debounce_clk_sel_out_mscbus;

// dp6 glitch filter bypass bus
input       [31:0] dp6_glitch_filter_bypass_out_mscbus;

// dp6 PES enable bus
input      [255:0] dp6_pes_en_out_mscbus;

// dp6 PES input enable bus
input       [31:0] dp6_pes_in_en_out_mscbus;

// dp6 PES safe value bus
input       [63:0] dp6_pes_safeval_out_mscbus;

// dp6 LVDS enable control bus
input       [31:0] dp6_lvds_en_ctrl_out_mscbus;

// dp6 input termination enable bus
input       [31:0] dp6_in_termination_en_out_mscbus;

// dp7 async input from pad bus
output      [31:0] dp7_async_in_from_pad_mscbus;

// dp7 gpio out to buf bus
input       [31:0] dp7_gpio_out_2_buf_mscbus;

// dp7 gpio out enable bus
input       [31:0] dp7_gpio_out_en_2_buf_mscbus;

// dp7 pinmux data to gpio bus
input       [31:0] dp7_pinmuxdata_2_gpio_mscbus;

// dp7 pinmux enable to gpio bus
input       [31:0] dp7_pinmuxen_2_gpio_mscbus;

// dp7 GP DATA IN out bus
output      [31:0] dp7_GP_DATA_IN_out_mscbus;

// dp7 data out to pinmux bus
output      [31:0] dp7_data_out_2_pinmux_mscbus;

// dp7 pinmux muxsel out bus
input      [159:0] dp7_pinmux_muxsel_out_mscbus;

// dp7 in function enable out bus
input     [1023:0] dp7_in_function_en_out_mscbus;

// dp7 analog mode select bus
input       [31:0] dp7_amsel_out_mscbus;

// dp7 drive strength 0 bus
input       [31:0] dp7_ds0_out_mscbus;

// dp7 drive strength 1 bus
input       [31:0] dp7_ds1_out_mscbus;

// dp7 slew control bus
input       [31:0] dp7_slew_out_mscbus;

// dp7 schmitt trigger bus
input       [31:0] dp7_schmitt_out_mscbus;

// dp7 mode 0 bus
input       [31:0] dp7_mode0_out_mscbus;

// dp7 mode 1 bus
input       [31:0] dp7_mode1_out_mscbus;

// dp7 input enable bus
input       [31:0] dp7_inena_out_mscbus;

// dp7 direction bus
input       [31:0] dp7_dir_out_mscbus;

// dp7 pull enable bus
input       [31:0] dp7_pull_en_out_mscbus;

// dp7 pull type bus
input       [31:0] dp7_pull_type_out_mscbus;

// dp7 glitch filter debounce clock select bus
input       [63:0] dp7_glitch_filter_debounce_clk_sel_out_mscbus;

// dp7 glitch filter bypass bus
input       [31:0] dp7_glitch_filter_bypass_out_mscbus;

// dp7 PES enable bus
input      [255:0] dp7_pes_en_out_mscbus;

// dp7 PES input enable bus
input       [31:0] dp7_pes_in_en_out_mscbus;

// dp7 PES safe value bus
input       [63:0] dp7_pes_safeval_out_mscbus;

// dp7 LVDS enable control bus
input       [31:0] dp7_lvds_en_ctrl_out_mscbus;

// dp7 input termination enable bus
input       [31:0] dp7_in_termination_en_out_mscbus;

// mp0 async input from pad bus
output      [31:0] mp0_async_in_from_pad_mscbus;

// mp0 gpio out to buf bus
input       [31:0] mp0_gpio_out_2_buf_mscbus;

// mp0 gpio out enable bus
input       [31:0] mp0_gpio_out_en_2_buf_mscbus;

// mp0 pinmux data to gpio bus
input       [31:0] mp0_pinmuxdata_2_gpio_mscbus;

// mp0 pinmux enable to gpio bus
input       [31:0] mp0_pinmuxen_2_gpio_mscbus;

// mp0 GP DATA IN out bus
output      [31:0] mp0_GP_DATA_IN_out_mscbus;

// mp0 data out to pinmux bus
output      [31:0] mp0_data_out_2_pinmux_mscbus;

// mp0 pinmux muxsel out bus
input      [159:0] mp0_pinmux_muxsel_out_mscbus;

// mp0 in function enable out bus
input     [1023:0] mp0_in_function_en_out_mscbus;

// mp0 analog mode select bus
input       [31:0] mp0_amsel_out_mscbus;

// mp0 drive strength 0 bus
input       [31:0] mp0_ds0_out_mscbus;

// mp0 drive strength 1 bus
input       [31:0] mp0_ds1_out_mscbus;

// mp0 slew control bus
input       [31:0] mp0_slew_out_mscbus;

// mp0 schmitt trigger bus
input       [31:0] mp0_schmitt_out_mscbus;

// mp0 mode 0 bus
input       [31:0] mp0_mode0_out_mscbus;

// mp0 mode 1 bus
input       [31:0] mp0_mode1_out_mscbus;

// mp0 input enable bus
input       [31:0] mp0_inena_out_mscbus;

// mp0 direction bus
input       [31:0] mp0_dir_out_mscbus;

// mp0 pull enable bus
input       [31:0] mp0_pull_en_out_mscbus;

// mp0 pull type bus
input       [31:0] mp0_pull_type_out_mscbus;

// mp0 glitch filter debounce clock select bus
input       [63:0] mp0_glitch_filter_debounce_clk_sel_out_mscbus;

// mp0 glitch filter bypass bus
input       [31:0] mp0_glitch_filter_bypass_out_mscbus;

// mp0 PES enable bus
input      [255:0] mp0_pes_en_out_mscbus;

// mp0 PES input enable bus
input       [31:0] mp0_pes_in_en_out_mscbus;

// mp0 PES safe value bus
input       [63:0] mp0_pes_safeval_out_mscbus;

// mp0 LVDS enable control bus
input       [31:0] mp0_lvds_en_ctrl_out_mscbus;

// mp0 input termination enable bus
input       [31:0] mp0_in_termination_en_out_mscbus;

// mp1 async input from pad bus
output      [31:0] mp1_async_in_from_pad_mscbus;

// mp1 gpio out to buf bus
input       [31:0] mp1_gpio_out_2_buf_mscbus;

// mp1 gpio out enable bus
input       [31:0] mp1_gpio_out_en_2_buf_mscbus;

// mp1 pinmux data to gpio bus
input       [31:0] mp1_pinmuxdata_2_gpio_mscbus;

// mp1 pinmux enable to gpio bus
input       [31:0] mp1_pinmuxen_2_gpio_mscbus;

// mp1 GP DATA IN out bus
output      [31:0] mp1_GP_DATA_IN_out_mscbus;

// mp1 data out to pinmux bus
output      [31:0] mp1_data_out_2_pinmux_mscbus;

// mp1 pinmux muxsel out bus
input      [159:0] mp1_pinmux_muxsel_out_mscbus;

// mp1 in function enable out bus
input     [1023:0] mp1_in_function_en_out_mscbus;

// mp1 analog mode select bus
input       [31:0] mp1_amsel_out_mscbus;

// mp1 drive strength 0 bus
input       [31:0] mp1_ds0_out_mscbus;

// mp1 drive strength 1 bus
input       [31:0] mp1_ds1_out_mscbus;

// mp1 slew control bus
input       [31:0] mp1_slew_out_mscbus;

// mp1 schmitt trigger bus
input       [31:0] mp1_schmitt_out_mscbus;

// mp1 mode 0 bus
input       [31:0] mp1_mode0_out_mscbus;

// mp1 mode 1 bus
input       [31:0] mp1_mode1_out_mscbus;

// mp1 input enable bus
input       [31:0] mp1_inena_out_mscbus;

// mp1 direction bus
input       [31:0] mp1_dir_out_mscbus;

// mp1 pull enable bus
input       [31:0] mp1_pull_en_out_mscbus;

// mp1 pull type bus
input       [31:0] mp1_pull_type_out_mscbus;

// mp1 glitch filter debounce clock select bus
input       [63:0] mp1_glitch_filter_debounce_clk_sel_out_mscbus;

// mp1 glitch filter bypass bus
input       [31:0] mp1_glitch_filter_bypass_out_mscbus;

// mp1 PES enable bus
input      [255:0] mp1_pes_en_out_mscbus;

// mp1 PES input enable bus
input       [31:0] mp1_pes_in_en_out_mscbus;

// mp1 PES safe value bus
input       [63:0] mp1_pes_safeval_out_mscbus;

// mp1 LVDS enable control bus
input       [31:0] mp1_lvds_en_ctrl_out_mscbus;

// mp1 input termination enable bus
input       [31:0] mp1_in_termination_en_out_mscbus;

// mp2 async input from pad bus
output      [31:0] mp2_async_in_from_pad_mscbus;

// mp2 gpio out to buf bus
input       [31:0] mp2_gpio_out_2_buf_mscbus;

// mp2 gpio out enable bus
input       [31:0] mp2_gpio_out_en_2_buf_mscbus;

// mp2 pinmux data to gpio bus
input       [31:0] mp2_pinmuxdata_2_gpio_mscbus;

// mp2 pinmux enable to gpio bus
input       [31:0] mp2_pinmuxen_2_gpio_mscbus;

// mp2 GP DATA IN out bus
output      [31:0] mp2_GP_DATA_IN_out_mscbus;

// mp2 data out to pinmux bus
output      [31:0] mp2_data_out_2_pinmux_mscbus;

// mp2 pinmux muxsel out bus
input      [159:0] mp2_pinmux_muxsel_out_mscbus;

// mp2 in function enable out bus
input     [1023:0] mp2_in_function_en_out_mscbus;

// mp2 analog mode select bus
input       [31:0] mp2_amsel_out_mscbus;

// mp2 drive strength 0 bus
input       [31:0] mp2_ds0_out_mscbus;

// mp2 drive strength 1 bus
input       [31:0] mp2_ds1_out_mscbus;

// mp2 slew control bus
input       [31:0] mp2_slew_out_mscbus;

// mp2 schmitt trigger bus
input       [31:0] mp2_schmitt_out_mscbus;

// mp2 mode 0 bus
input       [31:0] mp2_mode0_out_mscbus;

// mp2 mode 1 bus
input       [31:0] mp2_mode1_out_mscbus;

// mp2 input enable bus
input       [31:0] mp2_inena_out_mscbus;

// mp2 direction bus
input       [31:0] mp2_dir_out_mscbus;

// mp2 pull enable bus
input       [31:0] mp2_pull_en_out_mscbus;

// mp2 pull type bus
input       [31:0] mp2_pull_type_out_mscbus;

// mp2 glitch filter debounce clock select bus
input       [63:0] mp2_glitch_filter_debounce_clk_sel_out_mscbus;

// mp2 glitch filter bypass bus
input       [31:0] mp2_glitch_filter_bypass_out_mscbus;

// mp2 PES enable bus
input      [255:0] mp2_pes_en_out_mscbus;

// mp2 PES input enable bus
input       [31:0] mp2_pes_in_en_out_mscbus;

// mp2 PES safe value bus
input       [63:0] mp2_pes_safeval_out_mscbus;

// mp2 LVDS enable control bus
input       [31:0] mp2_lvds_en_ctrl_out_mscbus;

// mp2 input termination enable bus
input       [31:0] mp2_in_termination_en_out_mscbus;

// ap async input from pad bus
output      [31:0] ap_async_in_from_pad_mscbus;

// ap gpio out to buf bus
input       [31:0] ap_gpio_out_2_buf_mscbus;

// ap gpio out enable bus
input       [31:0] ap_gpio_out_en_2_buf_mscbus;

// ap pinmux data to gpio bus
input       [31:0] ap_pinmuxdata_2_gpio_mscbus;

// ap pinmux enable to gpio bus
input       [31:0] ap_pinmuxen_2_gpio_mscbus;

// ap GP DATA IN out bus
output      [31:0] ap_GP_DATA_IN_out_mscbus;

// ap data out to pinmux bus
output      [31:0] ap_data_out_2_pinmux_mscbus;

// ap pinmux muxsel out bus
input      [159:0] ap_pinmux_muxsel_out_mscbus;

// ap in function enable out bus
input     [1023:0] ap_in_function_en_out_mscbus;

// ap analog mode select bus
input       [31:0] ap_amsel_out_mscbus;

// ap drive strength 0 bus
input       [31:0] ap_ds0_out_mscbus;

// ap drive strength 1 bus
input       [31:0] ap_ds1_out_mscbus;

// ap slew control bus
input       [31:0] ap_slew_out_mscbus;

// ap schmitt trigger bus
input       [31:0] ap_schmitt_out_mscbus;

// ap mode 0 bus
input       [31:0] ap_mode0_out_mscbus;

// ap mode 1 bus
input       [31:0] ap_mode1_out_mscbus;

// ap input enable bus
input       [31:0] ap_inena_out_mscbus;

// ap direction bus
input       [31:0] ap_dir_out_mscbus;

// ap pull enable bus
input       [31:0] ap_pull_en_out_mscbus;

// ap pull type bus
input       [31:0] ap_pull_type_out_mscbus;

// ap glitch filter debounce clock select bus
input       [63:0] ap_glitch_filter_debounce_clk_sel_out_mscbus;

// ap glitch filter bypass bus
input       [31:0] ap_glitch_filter_bypass_out_mscbus;

// ap PES enable bus
input      [255:0] ap_pes_en_out_mscbus;

// ap PES input enable bus
input       [31:0] ap_pes_in_en_out_mscbus;

// ap PES safe value bus
input       [63:0] ap_pes_safeval_out_mscbus;

// ap LVDS enable control bus
input       [31:0] ap_lvds_en_ctrl_out_mscbus;

// ap input termination enable bus
input       [31:0] ap_in_termination_en_out_mscbus;

// DP0_0 input mux peripheral bus
input        [6:0] DP0_0_in_mux_peripheral_mscbus;

// DP0_1 input mux peripheral bus
input        [3:0] DP0_1_in_mux_peripheral_mscbus;

// DP0_1 output demux peripheral bus
output       [1:0] DP0_1_out_demux_peripheral_mscbus;

// DP0_2 input mux peripheral bus
input        [5:0] DP0_2_in_mux_peripheral_mscbus;

// DP0_3 input mux peripheral bus
input        [4:0] DP0_3_in_mux_peripheral_mscbus;

// DP0_3 output demux peripheral bus
output            DP0_3_out_demux_peripheral_mscbus;

// DP0_4 input mux peripheral bus
input        [5:0] DP0_4_in_mux_peripheral_mscbus;

// DP0_5 input mux peripheral bus
input        [4:0] DP0_5_in_mux_peripheral_mscbus;

// DP0_5 output demux peripheral bus
output            DP0_5_out_demux_peripheral_mscbus;

// DP0_6 input mux peripheral bus
input        [5:0] DP0_6_in_mux_peripheral_mscbus;

// DP0_7 input mux peripheral bus
input        [4:0] DP0_7_in_mux_peripheral_mscbus;

// DP0_7 output demux peripheral bus
output            DP0_7_out_demux_peripheral_mscbus;

// DP0_8 input mux peripheral bus
input        [4:0] DP0_8_in_mux_peripheral_mscbus;

// DP0_8 output demux peripheral bus
output            DP0_8_out_demux_peripheral_mscbus;

// DP0_9 input mux peripheral bus
input        [4:0] DP0_9_in_mux_peripheral_mscbus;

// DP0_9 output demux peripheral bus
output            DP0_9_out_demux_peripheral_mscbus;

// DP0_10 input mux peripheral bus
input        [4:0] DP0_10_in_mux_peripheral_mscbus;

// DP0_11 input mux peripheral bus
input        [4:0] DP0_11_in_mux_peripheral_mscbus;

// DP0_12 input mux peripheral bus
input        [4:0] DP0_12_in_mux_peripheral_mscbus;

// DP0_13 input mux peripheral bus
input        [4:0] DP0_13_in_mux_peripheral_mscbus;

// DP0_13 output demux peripheral bus
output            DP0_13_out_demux_peripheral_mscbus;

// DP0_14 input mux peripheral bus
input        [5:0] DP0_14_in_mux_peripheral_mscbus;

// DP0_14 output demux peripheral bus
output            DP0_14_out_demux_peripheral_mscbus;

// DP0_15 input mux peripheral bus
input        [5:0] DP0_15_in_mux_peripheral_mscbus;

// DP0_15 output demux peripheral bus
output            DP0_15_out_demux_peripheral_mscbus;

// DP0_16 input mux peripheral bus
input        [3:0] DP0_16_in_mux_peripheral_mscbus;

// DP0_16 output demux peripheral bus
output       [1:0] DP0_16_out_demux_peripheral_mscbus;

// DP0_17 input mux peripheral bus
input        [4:0] DP0_17_in_mux_peripheral_mscbus;

// DP0_17 output demux peripheral bus
output            DP0_17_out_demux_peripheral_mscbus;

// DP0_18 input mux peripheral bus
input        [4:0] DP0_18_in_mux_peripheral_mscbus;

// DP0_18 output demux peripheral bus
output            DP0_18_out_demux_peripheral_mscbus;

// DP0_19 input mux peripheral bus
input        [5:0] DP0_19_in_mux_peripheral_mscbus;

// DP0_20 input mux peripheral bus
input        [5:0] DP0_20_in_mux_peripheral_mscbus;

// DP0_21 input mux peripheral bus
input        [4:0] DP0_21_in_mux_peripheral_mscbus;

// DP0_21 output demux peripheral bus
output            DP0_21_out_demux_peripheral_mscbus;

// DP0_22 input mux peripheral bus
input        [3:0] DP0_22_in_mux_peripheral_mscbus;

// DP0_22 output demux peripheral bus
output       [1:0] DP0_22_out_demux_peripheral_mscbus;

// DP0_23 input mux peripheral bus
input        [3:0] DP0_23_in_mux_peripheral_mscbus;

// DP0_23 output demux peripheral bus
output       [1:0] DP0_23_out_demux_peripheral_mscbus;

// DP0_24 input mux peripheral bus
input        [3:0] DP0_24_in_mux_peripheral_mscbus;

// DP0_24 output demux peripheral bus
output       [1:0] DP0_24_out_demux_peripheral_mscbus;

// DP0_25 input mux peripheral bus
input        [4:0] DP0_25_in_mux_peripheral_mscbus;

// DP0_25 output demux peripheral bus
output            DP0_25_out_demux_peripheral_mscbus;

// DP0_26 input mux peripheral bus
input        [4:0] DP0_26_in_mux_peripheral_mscbus;

// DP0_26 output demux peripheral bus
output            DP0_26_out_demux_peripheral_mscbus;

// DP0_27 input mux peripheral bus
input        [4:0] DP0_27_in_mux_peripheral_mscbus;

// DP0_27 output demux peripheral bus
output            DP0_27_out_demux_peripheral_mscbus;

// DP0_28 input mux peripheral bus
input        [3:0] DP0_28_in_mux_peripheral_mscbus;

// DP0_28 output demux peripheral bus
output            DP0_28_out_demux_peripheral_mscbus;

// DP0_29 input mux peripheral bus
input        [2:0] DP0_29_in_mux_peripheral_mscbus;

// DP0_29 output demux peripheral bus
output       [1:0] DP0_29_out_demux_peripheral_mscbus;

// DP0_30 input mux peripheral bus
input        [2:0] DP0_30_in_mux_peripheral_mscbus;

// DP0_30 output demux peripheral bus
output       [1:0] DP0_30_out_demux_peripheral_mscbus;

// DP0_31 input mux peripheral bus
input        [3:0] DP0_31_in_mux_peripheral_mscbus;

// DP0_31 output demux peripheral bus
output            DP0_31_out_demux_peripheral_mscbus;

// DP1_0 input mux peripheral bus
input        [2:0] DP1_0_in_mux_peripheral_mscbus;

// DP1_0 output demux peripheral bus
output       [1:0] DP1_0_out_demux_peripheral_mscbus;

// DP1_1 input mux peripheral bus
input        [2:0] DP1_1_in_mux_peripheral_mscbus;

// DP1_1 output demux peripheral bus
output       [1:0] DP1_1_out_demux_peripheral_mscbus;

// DP1_2 input mux peripheral bus
input        [2:0] DP1_2_in_mux_peripheral_mscbus;

// DP1_2 output demux peripheral bus
output       [1:0] DP1_2_out_demux_peripheral_mscbus;

// DP1_3 input mux peripheral bus
input        [3:0] DP1_3_in_mux_peripheral_mscbus;

// DP1_3 output demux peripheral bus
output            DP1_3_out_demux_peripheral_mscbus;

// DP1_4 input mux peripheral bus
input        [3:0] DP1_4_in_mux_peripheral_mscbus;

// DP1_4 output demux peripheral bus
output            DP1_4_out_demux_peripheral_mscbus;

// DP1_5 input mux peripheral bus
input        [3:0] DP1_5_in_mux_peripheral_mscbus;

// DP1_5 output demux peripheral bus
output            DP1_5_out_demux_peripheral_mscbus;

// DP1_6 input mux peripheral bus
input        [2:0] DP1_6_in_mux_peripheral_mscbus;

// DP1_6 output demux peripheral bus
output       [1:0] DP1_6_out_demux_peripheral_mscbus;

// DP1_7 input mux peripheral bus
input        [3:0] DP1_7_in_mux_peripheral_mscbus;

// DP1_7 output demux peripheral bus
output            DP1_7_out_demux_peripheral_mscbus;

// DP1_8 input mux peripheral bus
input        [2:0] DP1_8_in_mux_peripheral_mscbus;

// DP1_8 output demux peripheral bus
output            DP1_8_out_demux_peripheral_mscbus;

// DP1_9 input mux peripheral bus
input        [2:0] DP1_9_in_mux_peripheral_mscbus;

// DP1_9 output demux peripheral bus
output            DP1_9_out_demux_peripheral_mscbus;

// DP1_10 input mux peripheral bus
input        [1:0] DP1_10_in_mux_peripheral_mscbus;

// DP1_10 output demux peripheral bus
output       [1:0] DP1_10_out_demux_peripheral_mscbus;

// DP1_11 input mux peripheral bus
input        [1:0] DP1_11_in_mux_peripheral_mscbus;

// DP1_11 output demux peripheral bus
output       [1:0] DP1_11_out_demux_peripheral_mscbus;

// DP1_12 input mux peripheral bus
input        [1:0] DP1_12_in_mux_peripheral_mscbus;

// DP1_12 output demux peripheral bus
output            DP1_12_out_demux_peripheral_mscbus;

// DP1_13 input mux peripheral bus
input        [3:0] DP1_13_in_mux_peripheral_mscbus;

// DP1_13 output demux peripheral bus
output            DP1_13_out_demux_peripheral_mscbus;

// DP1_14 input mux peripheral bus
input        [1:0] DP1_14_in_mux_peripheral_mscbus;

// DP1_14 output demux peripheral bus
output       [2:0] DP1_14_out_demux_peripheral_mscbus;

// DP1_15 input mux peripheral bus
input        [3:0] DP1_15_in_mux_peripheral_mscbus;

// DP1_15 output demux peripheral bus
output            DP1_15_out_demux_peripheral_mscbus;

// DP1_16 input mux peripheral bus
input        [2:0] DP1_16_in_mux_peripheral_mscbus;

// DP1_16 output demux peripheral bus
output       [1:0] DP1_16_out_demux_peripheral_mscbus;

// DP1_17 input mux peripheral bus
input        [2:0] DP1_17_in_mux_peripheral_mscbus;

// DP1_17 output demux peripheral bus
output       [1:0] DP1_17_out_demux_peripheral_mscbus;

// DP1_18 input mux peripheral bus
input        [2:0] DP1_18_in_mux_peripheral_mscbus;

// DP1_18 output demux peripheral bus
output       [1:0] DP1_18_out_demux_peripheral_mscbus;

// DP1_19 input mux peripheral bus
input        [3:0] DP1_19_in_mux_peripheral_mscbus;

// DP1_19 output demux peripheral bus
output            DP1_19_out_demux_peripheral_mscbus;

// DP1_20 input mux peripheral bus
input        [2:0] DP1_20_in_mux_peripheral_mscbus;

// DP1_20 output demux peripheral bus
output       [1:0] DP1_20_out_demux_peripheral_mscbus;

// DP1_21 input mux peripheral bus
input        [3:0] DP1_21_in_mux_peripheral_mscbus;

// DP1_21 output demux peripheral bus
output            DP1_21_out_demux_peripheral_mscbus;

// DP1_22 input mux peripheral bus
input        [3:0] DP1_22_in_mux_peripheral_mscbus;

// DP1_22 output demux peripheral bus
output            DP1_22_out_demux_peripheral_mscbus;

// DP1_23 input mux peripheral bus
input        [2:0] DP1_23_in_mux_peripheral_mscbus;

// DP1_23 output demux peripheral bus
output            DP1_23_out_demux_peripheral_mscbus;

// DP1_24 input mux peripheral bus
input        [2:0] DP1_24_in_mux_peripheral_mscbus;

// DP1_24 output demux peripheral bus
output            DP1_24_out_demux_peripheral_mscbus;

// DP1_25 input mux peripheral bus
input        [4:0] DP1_25_in_mux_peripheral_mscbus;

// DP1_26 input mux peripheral bus
input        [4:0] DP1_26_in_mux_peripheral_mscbus;

// DP1_27 input mux peripheral bus
input        [4:0] DP1_27_in_mux_peripheral_mscbus;

// DP1_28 input mux peripheral bus
input        [3:0] DP1_28_in_mux_peripheral_mscbus;

// DP1_28 output demux peripheral bus
output            DP1_28_out_demux_peripheral_mscbus;

// DP1_29 input mux peripheral bus
input        [3:0] DP1_29_in_mux_peripheral_mscbus;

// DP1_29 output demux peripheral bus
output            DP1_29_out_demux_peripheral_mscbus;

// DP1_30 input mux peripheral bus
input        [3:0] DP1_30_in_mux_peripheral_mscbus;

// DP1_30 output demux peripheral bus
output            DP1_30_out_demux_peripheral_mscbus;

// DP1_31 input mux peripheral bus
input        [2:0] DP1_31_in_mux_peripheral_mscbus;

// DP1_31 output demux peripheral bus
output       [1:0] DP1_31_out_demux_peripheral_mscbus;

// DP2_0 input mux peripheral bus
input        [3:0] DP2_0_in_mux_peripheral_mscbus;

// DP2_0 output demux peripheral bus
output            DP2_0_out_demux_peripheral_mscbus;

// DP2_1 input mux peripheral bus
input        [3:0] DP2_1_in_mux_peripheral_mscbus;

// DP2_2 input mux peripheral bus
input        [3:0] DP2_2_in_mux_peripheral_mscbus;

// DP2_2 output demux peripheral bus
output            DP2_2_out_demux_peripheral_mscbus;

// DP2_3 input mux peripheral bus
input        [3:0] DP2_3_in_mux_peripheral_mscbus;

// DP2_3 output demux peripheral bus
output            DP2_3_out_demux_peripheral_mscbus;

// DP2_4 input mux peripheral bus
input        [3:0] DP2_4_in_mux_peripheral_mscbus;

// DP2_5 input mux peripheral bus
input        [3:0] DP2_5_in_mux_peripheral_mscbus;

// DP2_6 input mux peripheral bus
input        [2:0] DP2_6_in_mux_peripheral_mscbus;

// DP2_6 output demux peripheral bus
output            DP2_6_out_demux_peripheral_mscbus;

// DP2_7 input mux peripheral bus
input        [3:0] DP2_7_in_mux_peripheral_mscbus;

// DP2_8 input mux peripheral bus
input        [3:0] DP2_8_in_mux_peripheral_mscbus;

// DP2_9 input mux peripheral bus
input        [3:0] DP2_9_in_mux_peripheral_mscbus;

// DP2_10 input mux peripheral bus
input        [3:0] DP2_10_in_mux_peripheral_mscbus;

// DP2_11 input mux peripheral bus
input        [2:0] DP2_11_in_mux_peripheral_mscbus;

// DP2_12 input mux peripheral bus
input        [3:0] DP2_12_in_mux_peripheral_mscbus;

// DP2_12 output demux peripheral bus
output            DP2_12_out_demux_peripheral_mscbus;

// DP2_13 input mux peripheral bus
input        [2:0] DP2_13_in_mux_peripheral_mscbus;

// DP2_13 output demux peripheral bus
output            DP2_13_out_demux_peripheral_mscbus;

// DP2_14 input mux peripheral bus
input        [3:0] DP2_14_in_mux_peripheral_mscbus;

// DP2_15 input mux peripheral bus
input        [2:0] DP2_15_in_mux_peripheral_mscbus;

// DP2_15 output demux peripheral bus
output            DP2_15_out_demux_peripheral_mscbus;

// DP2_16 input mux peripheral bus
input        [2:0] DP2_16_in_mux_peripheral_mscbus;

// DP2_16 output demux peripheral bus
output            DP2_16_out_demux_peripheral_mscbus;

// DP2_17 input mux peripheral bus
input        [2:0] DP2_17_in_mux_peripheral_mscbus;

// DP2_17 output demux peripheral bus
output            DP2_17_out_demux_peripheral_mscbus;

// DP2_18 input mux peripheral bus
input        [3:0] DP2_18_in_mux_peripheral_mscbus;

// DP2_19 input mux peripheral bus
input        [3:0] DP2_19_in_mux_peripheral_mscbus;

// DP2_20 input mux peripheral bus
input        [2:0] DP2_20_in_mux_peripheral_mscbus;

// DP2_20 output demux peripheral bus
output            DP2_20_out_demux_peripheral_mscbus;

// DP2_21 input mux peripheral bus
input        [5:0] DP2_21_in_mux_peripheral_mscbus;

// DP2_22 input mux peripheral bus
input        [4:0] DP2_22_in_mux_peripheral_mscbus;

// DP2_22 output demux peripheral bus
output            DP2_22_out_demux_peripheral_mscbus;

// DP2_23 input mux peripheral bus
input        [5:0] DP2_23_in_mux_peripheral_mscbus;

// DP2_23 output demux peripheral bus
output            DP2_23_out_demux_peripheral_mscbus;

// DP2_24 input mux peripheral bus
input        [4:0] DP2_24_in_mux_peripheral_mscbus;

// DP2_24 output demux peripheral bus
output       [1:0] DP2_24_out_demux_peripheral_mscbus;

// DP2_25 input mux peripheral bus
input        [5:0] DP2_25_in_mux_peripheral_mscbus;

// DP2_26 input mux peripheral bus
input        [3:0] DP2_26_in_mux_peripheral_mscbus;

// DP2_26 output demux peripheral bus
output       [1:0] DP2_26_out_demux_peripheral_mscbus;

// DP2_27 input mux peripheral bus
input        [4:0] DP2_27_in_mux_peripheral_mscbus;

// DP2_27 output demux peripheral bus
output            DP2_27_out_demux_peripheral_mscbus;

// DP2_28 input mux peripheral bus
input        [2:0] DP2_28_in_mux_peripheral_mscbus;

// DP2_28 output demux peripheral bus
output       [2:0] DP2_28_out_demux_peripheral_mscbus;

// DP2_29 input mux peripheral bus
input        [4:0] DP2_29_in_mux_peripheral_mscbus;

// DP2_29 output demux peripheral bus
output            DP2_29_out_demux_peripheral_mscbus;

// DP2_30 input mux peripheral bus
input        [3:0] DP2_30_in_mux_peripheral_mscbus;

// DP2_30 output demux peripheral bus
output       [1:0] DP2_30_out_demux_peripheral_mscbus;

// DP2_31 input mux peripheral bus
input        [4:0] DP2_31_in_mux_peripheral_mscbus;

// DP2_31 output demux peripheral bus
output            DP2_31_out_demux_peripheral_mscbus;

// DP3_0 input mux peripheral bus
input        [3:0] DP3_0_in_mux_peripheral_mscbus;

// DP3_0 output demux peripheral bus
output       [1:0] DP3_0_out_demux_peripheral_mscbus;

// DP3_1 input mux peripheral bus
input        [3:0] DP3_1_in_mux_peripheral_mscbus;

// DP3_1 output demux peripheral bus
output       [1:0] DP3_1_out_demux_peripheral_mscbus;

// DP3_2 input mux peripheral bus
input        [4:0] DP3_2_in_mux_peripheral_mscbus;

// DP3_2 output demux peripheral bus
output            DP3_2_out_demux_peripheral_mscbus;

// DP3_3 input mux peripheral bus
input        [2:0] DP3_3_in_mux_peripheral_mscbus;

// DP3_3 output demux peripheral bus
output       [2:0] DP3_3_out_demux_peripheral_mscbus;

// DP3_4 input mux peripheral bus
input        [4:0] DP3_4_in_mux_peripheral_mscbus;

// DP3_4 output demux peripheral bus
output            DP3_4_out_demux_peripheral_mscbus;

// DP3_5 input mux peripheral bus
input        [3:0] DP3_5_in_mux_peripheral_mscbus;

// DP3_5 output demux peripheral bus
output            DP3_5_out_demux_peripheral_mscbus;

// DP3_6 input mux peripheral bus
input        [3:0] DP3_6_in_mux_peripheral_mscbus;

// DP3_6 output demux peripheral bus
output            DP3_6_out_demux_peripheral_mscbus;

// DP3_7 input mux peripheral bus
input        [3:0] DP3_7_in_mux_peripheral_mscbus;

// DP3_7 output demux peripheral bus
output            DP3_7_out_demux_peripheral_mscbus;

// DP3_8 input mux peripheral bus
input        [4:0] DP3_8_in_mux_peripheral_mscbus;

// DP3_8 output demux peripheral bus
output            DP3_8_out_demux_peripheral_mscbus;

// DP3_9 input mux peripheral bus
input        [3:0] DP3_9_in_mux_peripheral_mscbus;

// DP3_9 output demux peripheral bus
output       [1:0] DP3_9_out_demux_peripheral_mscbus;

// DP3_10 input mux peripheral bus
input        [2:0] DP3_10_in_mux_peripheral_mscbus;

// DP3_10 output demux peripheral bus
output       [2:0] DP3_10_out_demux_peripheral_mscbus;

// DP3_11 input mux peripheral bus
input        [3:0] DP3_11_in_mux_peripheral_mscbus;

// DP3_11 output demux peripheral bus
output       [1:0] DP3_11_out_demux_peripheral_mscbus;

// DP3_12 input mux peripheral bus
input        [5:0] DP3_12_in_mux_peripheral_mscbus;

// DP3_13 input mux peripheral bus
input        [3:0] DP3_13_in_mux_peripheral_mscbus;

// DP3_13 output demux peripheral bus
output       [1:0] DP3_13_out_demux_peripheral_mscbus;

// DP3_14 input mux peripheral bus
input        [5:0] DP3_14_in_mux_peripheral_mscbus;

// DP3_15 input mux peripheral bus
input        [4:0] DP3_15_in_mux_peripheral_mscbus;

// DP3_15 output demux peripheral bus
output            DP3_15_out_demux_peripheral_mscbus;

// DP3_16 input mux peripheral bus
input        [4:0] DP3_16_in_mux_peripheral_mscbus;

// DP3_16 output demux peripheral bus
output            DP3_16_out_demux_peripheral_mscbus;

// DP3_17 input mux peripheral bus
input        [3:0] DP3_17_in_mux_peripheral_mscbus;

// DP3_17 output demux peripheral bus
output       [1:0] DP3_17_out_demux_peripheral_mscbus;

// DP3_18 input mux peripheral bus
input        [5:0] DP3_18_in_mux_peripheral_mscbus;

// DP3_19 input mux peripheral bus
input        [5:0] DP3_19_in_mux_peripheral_mscbus;

// DP3_20 input mux peripheral bus
input        [5:0] DP3_20_in_mux_peripheral_mscbus;

// DP3_21 input mux peripheral bus
input        [6:0] DP3_21_in_mux_peripheral_mscbus;

// DP3_22 input mux peripheral bus
input        [6:0] DP3_22_in_mux_peripheral_mscbus;

// DP3_23 input mux peripheral bus
input        [6:0] DP3_23_in_mux_peripheral_mscbus;

// DP3_24 input mux peripheral bus
input        [4:0] DP3_24_in_mux_peripheral_mscbus;

// DP3_24 output demux peripheral bus
output       [1:0] DP3_24_out_demux_peripheral_mscbus;

// DP3_25 input mux peripheral bus
input        [5:0] DP3_25_in_mux_peripheral_mscbus;

// DP3_25 output demux peripheral bus
output            DP3_25_out_demux_peripheral_mscbus;

// DP3_26 input mux peripheral bus
input        [4:0] DP3_26_in_mux_peripheral_mscbus;

// DP3_26 output demux peripheral bus
output       [1:0] DP3_26_out_demux_peripheral_mscbus;

// DP3_27 input mux peripheral bus
input        [4:0] DP3_27_in_mux_peripheral_mscbus;

// DP3_27 output demux peripheral bus
output       [1:0] DP3_27_out_demux_peripheral_mscbus;

// DP3_28 input mux peripheral bus
input        [4:0] DP3_28_in_mux_peripheral_mscbus;

// DP3_28 output demux peripheral bus
output       [1:0] DP3_28_out_demux_peripheral_mscbus;

// DP3_29 input mux peripheral bus
input        [4:0] DP3_29_in_mux_peripheral_mscbus;

// DP3_30 input mux peripheral bus
input        [4:0] DP3_30_in_mux_peripheral_mscbus;

// DP3_30 output demux peripheral bus
output            DP3_30_out_demux_peripheral_mscbus;

// DP3_31 input mux peripheral bus
input        [2:0] DP3_31_in_mux_peripheral_mscbus;

// DP3_31 output demux peripheral bus
output       [2:0] DP3_31_out_demux_peripheral_mscbus;

// DP4_0 input mux peripheral bus
input        [3:0] DP4_0_in_mux_peripheral_mscbus;

// DP4_0 output demux peripheral bus
output            DP4_0_out_demux_peripheral_mscbus;

// DP4_1 input mux peripheral bus
input        [2:0] DP4_1_in_mux_peripheral_mscbus;

// DP4_1 output demux peripheral bus
output       [1:0] DP4_1_out_demux_peripheral_mscbus;

// DP4_2 input mux peripheral bus
input        [3:0] DP4_2_in_mux_peripheral_mscbus;

// DP4_2 output demux peripheral bus
output            DP4_2_out_demux_peripheral_mscbus;

// DP4_3 input mux peripheral bus
input        [3:0] DP4_3_in_mux_peripheral_mscbus;

// DP4_3 output demux peripheral bus
output            DP4_3_out_demux_peripheral_mscbus;

// DP4_4 input mux peripheral bus
input        [2:0] DP4_4_in_mux_peripheral_mscbus;

// DP4_4 output demux peripheral bus
output       [1:0] DP4_4_out_demux_peripheral_mscbus;

// DP4_5 input mux peripheral bus
input        [4:0] DP4_5_in_mux_peripheral_mscbus;

// DP4_6 input mux peripheral bus
input        [5:0] DP4_6_in_mux_peripheral_mscbus;

// DP4_6 output demux peripheral bus
output       [1:0] DP4_6_out_demux_peripheral_mscbus;

// DP4_7 input mux peripheral bus
input        [5:0] DP4_7_in_mux_peripheral_mscbus;

// DP4_7 output demux peripheral bus
output            DP4_7_out_demux_peripheral_mscbus;

// DP4_8 input mux peripheral bus
input        [6:0] DP4_8_in_mux_peripheral_mscbus;

// DP4_9 input mux peripheral bus
input        [4:0] DP4_9_in_mux_peripheral_mscbus;

// DP4_9 output demux peripheral bus
output       [1:0] DP4_9_out_demux_peripheral_mscbus;

// DP4_10 input mux peripheral bus
input        [4:0] DP4_10_in_mux_peripheral_mscbus;

// DP4_10 output demux peripheral bus
output       [1:0] DP4_10_out_demux_peripheral_mscbus;

// DP4_11 input mux peripheral bus
input        [5:0] DP4_11_in_mux_peripheral_mscbus;

// DP4_11 output demux peripheral bus
output            DP4_11_out_demux_peripheral_mscbus;

// DP4_12 input mux peripheral bus
input        [4:0] DP4_12_in_mux_peripheral_mscbus;

// DP4_12 output demux peripheral bus
output       [1:0] DP4_12_out_demux_peripheral_mscbus;

// DP4_13 input mux peripheral bus
input        [4:0] DP4_13_in_mux_peripheral_mscbus;

// DP4_13 output demux peripheral bus
output       [1:0] DP4_13_out_demux_peripheral_mscbus;

// DP4_14 input mux peripheral bus
input        [3:0] DP4_14_in_mux_peripheral_mscbus;

// DP4_14 output demux peripheral bus
output            DP4_14_out_demux_peripheral_mscbus;

// DP4_15 input mux peripheral bus
input        [3:0] DP4_15_in_mux_peripheral_mscbus;

// DP4_15 output demux peripheral bus
output       [2:0] DP4_15_out_demux_peripheral_mscbus;

// DP4_16 input mux peripheral bus
input        [3:0] DP4_16_in_mux_peripheral_mscbus;

// DP4_16 output demux peripheral bus
output       [2:0] DP4_16_out_demux_peripheral_mscbus;

// DP4_17 input mux peripheral bus
input        [3:0] DP4_17_in_mux_peripheral_mscbus;

// DP4_17 output demux peripheral bus
output       [2:0] DP4_17_out_demux_peripheral_mscbus;

// DP4_18 input mux peripheral bus
input        [1:0] DP4_18_in_mux_peripheral_mscbus;

// DP4_18 output demux peripheral bus
output       [1:0] DP4_18_out_demux_peripheral_mscbus;

// DP4_19 input mux peripheral bus
input        [2:0] DP4_19_in_mux_peripheral_mscbus;

// DP4_20 input mux peripheral bus
input        [5:0] DP4_20_in_mux_peripheral_mscbus;

// DP4_21 input mux peripheral bus
input        [5:0] DP4_21_in_mux_peripheral_mscbus;

// DP4_22 input mux peripheral bus
input        [4:0] DP4_22_in_mux_peripheral_mscbus;

// DP4_22 output demux peripheral bus
output            DP4_22_out_demux_peripheral_mscbus;

// DP4_23 input mux peripheral bus
input        [4:0] DP4_23_in_mux_peripheral_mscbus;

// DP4_24 input mux peripheral bus
input        [4:0] DP4_24_in_mux_peripheral_mscbus;

// DP4_25 input mux peripheral bus
input        [2:0] DP4_25_in_mux_peripheral_mscbus;

// DP4_25 output demux peripheral bus
output            DP4_25_out_demux_peripheral_mscbus;

// DP4_26 input mux peripheral bus
input        [3:0] DP4_26_in_mux_peripheral_mscbus;

// DP4_27 input mux peripheral bus
input        [3:0] DP4_27_in_mux_peripheral_mscbus;

// DP4_27 output demux peripheral bus
output            DP4_27_out_demux_peripheral_mscbus;

// DP4_28 input mux peripheral bus
input        [4:0] DP4_28_in_mux_peripheral_mscbus;

// DP4_28 output demux peripheral bus
output            DP4_28_out_demux_peripheral_mscbus;

// DP4_29 input mux peripheral bus
input        [2:0] DP4_29_in_mux_peripheral_mscbus;

// DP4_29 output demux peripheral bus
output       [1:0] DP4_29_out_demux_peripheral_mscbus;

// DP4_30 input mux peripheral bus
input        [3:0] DP4_30_in_mux_peripheral_mscbus;

// DP4_30 output demux peripheral bus
output            DP4_30_out_demux_peripheral_mscbus;

// DP4_31 input mux peripheral bus
input        [2:0] DP4_31_in_mux_peripheral_mscbus;

// DP4_31 output demux peripheral bus
output       [1:0] DP4_31_out_demux_peripheral_mscbus;

// DP5_0 input mux peripheral bus
input        [6:0] DP5_0_in_mux_peripheral_mscbus;

// DP5_1 input mux peripheral bus
input        [4:0] DP5_1_in_mux_peripheral_mscbus;

// DP5_1 output demux peripheral bus
output            DP5_1_out_demux_peripheral_mscbus;

// DP5_2 input mux peripheral bus
input        [4:0] DP5_2_in_mux_peripheral_mscbus;

// DP5_2 output demux peripheral bus
output            DP5_2_out_demux_peripheral_mscbus;

// DP5_3 input mux peripheral bus
input        [4:0] DP5_3_in_mux_peripheral_mscbus;

// DP5_3 output demux peripheral bus
output            DP5_3_out_demux_peripheral_mscbus;

// DP5_4 input mux peripheral bus
input        [4:0] DP5_4_in_mux_peripheral_mscbus;

// DP5_4 output demux peripheral bus
output       [1:0] DP5_4_out_demux_peripheral_mscbus;

// DP5_5 input mux peripheral bus
input        [4:0] DP5_5_in_mux_peripheral_mscbus;

// DP5_5 output demux peripheral bus
output       [1:0] DP5_5_out_demux_peripheral_mscbus;

// DP5_6 input mux peripheral bus
input        [6:0] DP5_6_in_mux_peripheral_mscbus;

// DP5_6 output demux peripheral bus
output            DP5_6_out_demux_peripheral_mscbus;

// DP5_7 input mux peripheral bus
input        [6:0] DP5_7_in_mux_peripheral_mscbus;

// DP5_8 input mux peripheral bus
input        [5:0] DP5_8_in_mux_peripheral_mscbus;

// DP5_8 output demux peripheral bus
output            DP5_8_out_demux_peripheral_mscbus;

// DP5_9 input mux peripheral bus
input        [2:0] DP5_9_in_mux_peripheral_mscbus;

// DP5_9 output demux peripheral bus
output       [3:0] DP5_9_out_demux_peripheral_mscbus;

// DP5_10 input mux peripheral bus
input        [4:0] DP5_10_in_mux_peripheral_mscbus;

// DP5_10 output demux peripheral bus
output       [1:0] DP5_10_out_demux_peripheral_mscbus;

// DP5_11 input mux peripheral bus
input        [3:0] DP5_11_in_mux_peripheral_mscbus;

// DP5_11 output demux peripheral bus
output       [2:0] DP5_11_out_demux_peripheral_mscbus;

// DP5_12 input mux peripheral bus
input        [4:0] DP5_12_in_mux_peripheral_mscbus;

// DP5_12 output demux peripheral bus
output       [1:0] DP5_12_out_demux_peripheral_mscbus;

// DP5_13 input mux peripheral bus
input        [4:0] DP5_13_in_mux_peripheral_mscbus;

// DP5_13 output demux peripheral bus
output       [1:0] DP5_13_out_demux_peripheral_mscbus;

// DP5_14 input mux peripheral bus
input        [5:0] DP5_14_in_mux_peripheral_mscbus;

// DP5_15 input mux peripheral bus
input        [4:0] DP5_15_in_mux_peripheral_mscbus;

// DP5_15 output demux peripheral bus
output            DP5_15_out_demux_peripheral_mscbus;

// DP5_16 input mux peripheral bus
input        [4:0] DP5_16_in_mux_peripheral_mscbus;

// DP5_16 output demux peripheral bus
output            DP5_16_out_demux_peripheral_mscbus;

// DP5_17 input mux peripheral bus
input        [4:0] DP5_17_in_mux_peripheral_mscbus;

// DP5_17 output demux peripheral bus
output            DP5_17_out_demux_peripheral_mscbus;

// DP5_18 input mux peripheral bus
input        [4:0] DP5_18_in_mux_peripheral_mscbus;

// DP5_19 input mux peripheral bus
input        [3:0] DP5_19_in_mux_peripheral_mscbus;

// DP5_19 output demux peripheral bus
output            DP5_19_out_demux_peripheral_mscbus;

// DP5_20 input mux peripheral bus
input        [5:0] DP5_20_in_mux_peripheral_mscbus;

// DP5_21 input mux peripheral bus
input        [4:0] DP5_21_in_mux_peripheral_mscbus;

// DP5_21 output demux peripheral bus
output            DP5_21_out_demux_peripheral_mscbus;

// DP5_22 input mux peripheral bus
input        [3:0] DP5_22_in_mux_peripheral_mscbus;

// DP5_22 output demux peripheral bus
output       [1:0] DP5_22_out_demux_peripheral_mscbus;

// DP5_23 input mux peripheral bus
input        [4:0] DP5_23_in_mux_peripheral_mscbus;

// DP5_23 output demux peripheral bus
output            DP5_23_out_demux_peripheral_mscbus;

// DP5_24 input mux peripheral bus
input        [4:0] DP5_24_in_mux_peripheral_mscbus;

// DP5_24 output demux peripheral bus
output            DP5_24_out_demux_peripheral_mscbus;

// DP5_25 input mux peripheral bus
input        [3:0] DP5_25_in_mux_peripheral_mscbus;

// DP5_25 output demux peripheral bus
output            DP5_25_out_demux_peripheral_mscbus;

// DP5_26 input mux peripheral bus
input        [5:0] DP5_26_in_mux_peripheral_mscbus;

// DP5_26 output demux peripheral bus
output            DP5_26_out_demux_peripheral_mscbus;

// DP5_27 input mux peripheral bus
input        [7:0] DP5_27_in_mux_peripheral_mscbus;

// DP5_28 input mux peripheral bus
input        [5:0] DP5_28_in_mux_peripheral_mscbus;

// DP5_28 output demux peripheral bus
output       [1:0] DP5_28_out_demux_peripheral_mscbus;

// DP5_29 input mux peripheral bus
input        [6:0] DP5_29_in_mux_peripheral_mscbus;

// DP5_29 output demux peripheral bus
output            DP5_29_out_demux_peripheral_mscbus;

// DP5_30 input mux peripheral bus
input        [4:0] DP5_30_in_mux_peripheral_mscbus;

// DP5_30 output demux peripheral bus
output       [2:0] DP5_30_out_demux_peripheral_mscbus;

// DP5_31 input mux peripheral bus
input        [6:0] DP5_31_in_mux_peripheral_mscbus;

// DP5_31 output demux peripheral bus
output            DP5_31_out_demux_peripheral_mscbus;

// DP6_0 input mux peripheral bus
input        [4:0] DP6_0_in_mux_peripheral_mscbus;

// DP6_0 output demux peripheral bus
output       [2:0] DP6_0_out_demux_peripheral_mscbus;

// DP6_1 input mux peripheral bus
input        [4:0] DP6_1_in_mux_peripheral_mscbus;

// DP6_1 output demux peripheral bus
output       [1:0] DP6_1_out_demux_peripheral_mscbus;

// DP6_2 input mux peripheral bus
input        [4:0] DP6_2_in_mux_peripheral_mscbus;

// DP6_2 output demux peripheral bus
output       [2:0] DP6_2_out_demux_peripheral_mscbus;

// DP6_3 input mux peripheral bus
input        [6:0] DP6_3_in_mux_peripheral_mscbus;

// DP6_3 output demux peripheral bus
output            DP6_3_out_demux_peripheral_mscbus;

// DP6_4 input mux peripheral bus
input        [4:0] DP6_4_in_mux_peripheral_mscbus;

// DP6_4 output demux peripheral bus
output       [1:0] DP6_4_out_demux_peripheral_mscbus;

// DP6_5 input mux peripheral bus
input        [4:0] DP6_5_in_mux_peripheral_mscbus;

// DP6_5 output demux peripheral bus
output       [1:0] DP6_5_out_demux_peripheral_mscbus;

// DP6_6 input mux peripheral bus
input        [5:0] DP6_6_in_mux_peripheral_mscbus;

// DP6_6 output demux peripheral bus
output            DP6_6_out_demux_peripheral_mscbus;

// DP6_7 input mux peripheral bus
input        [5:0] DP6_7_in_mux_peripheral_mscbus;

// DP6_7 output demux peripheral bus
output            DP6_7_out_demux_peripheral_mscbus;

// DP6_8 input mux peripheral bus
input        [3:0] DP6_8_in_mux_peripheral_mscbus;

// DP6_8 output demux peripheral bus
output       [1:0] DP6_8_out_demux_peripheral_mscbus;

// DP6_9 input mux peripheral bus
input        [4:0] DP6_9_in_mux_peripheral_mscbus;

// DP6_9 output demux peripheral bus
output            DP6_9_out_demux_peripheral_mscbus;

// DP6_10 input mux peripheral bus
input        [4:0] DP6_10_in_mux_peripheral_mscbus;

// DP6_10 output demux peripheral bus
output            DP6_10_out_demux_peripheral_mscbus;

// DP6_11 input mux peripheral bus
input        [5:0] DP6_11_in_mux_peripheral_mscbus;

// DP6_12 input mux peripheral bus
input        [5:0] DP6_12_in_mux_peripheral_mscbus;

// DP6_12 output demux peripheral bus
output            DP6_12_out_demux_peripheral_mscbus;

// DP6_13 input mux peripheral bus
input        [5:0] DP6_13_in_mux_peripheral_mscbus;

// DP6_13 output demux peripheral bus
output       [1:0] DP6_13_out_demux_peripheral_mscbus;

// DP6_14 input mux peripheral bus
input        [5:0] DP6_14_in_mux_peripheral_mscbus;

// DP6_14 output demux peripheral bus
output            DP6_14_out_demux_peripheral_mscbus;

// DP6_15 input mux peripheral bus
input        [4:0] DP6_15_in_mux_peripheral_mscbus;

// DP6_15 output demux peripheral bus
output       [1:0] DP6_15_out_demux_peripheral_mscbus;

// DP6_16 input mux peripheral bus
input        [5:0] DP6_16_in_mux_peripheral_mscbus;

// DP6_16 output demux peripheral bus
output            DP6_16_out_demux_peripheral_mscbus;

// DP6_17 input mux peripheral bus
input        [6:0] DP6_17_in_mux_peripheral_mscbus;

// DP6_18 input mux peripheral bus
input        [6:0] DP6_18_in_mux_peripheral_mscbus;

// DP6_18 output demux peripheral bus
output            DP6_18_out_demux_peripheral_mscbus;

// DP6_19 input mux peripheral bus
input        [4:0] DP6_19_in_mux_peripheral_mscbus;

// DP6_19 output demux peripheral bus
output       [1:0] DP6_19_out_demux_peripheral_mscbus;

// DP6_20 input mux peripheral bus
input        [6:0] DP6_20_in_mux_peripheral_mscbus;

// DP6_21 input mux peripheral bus
input        [3:0] DP6_21_in_mux_peripheral_mscbus;

// DP6_21 output demux peripheral bus
output       [2:0] DP6_21_out_demux_peripheral_mscbus;

// DP6_22 input mux peripheral bus
input        [4:0] DP6_22_in_mux_peripheral_mscbus;

// DP6_22 output demux peripheral bus
output       [1:0] DP6_22_out_demux_peripheral_mscbus;

// DP6_23 input mux peripheral bus
input        [5:0] DP6_23_in_mux_peripheral_mscbus;

// DP6_23 output demux peripheral bus
output            DP6_23_out_demux_peripheral_mscbus;

// DP6_24 input mux peripheral bus
input        [5:0] DP6_24_in_mux_peripheral_mscbus;

// DP6_24 output demux peripheral bus
output            DP6_24_out_demux_peripheral_mscbus;

// DP6_25 input mux peripheral bus
input        [4:0] DP6_25_in_mux_peripheral_mscbus;

// DP6_25 output demux peripheral bus
output       [1:0] DP6_25_out_demux_peripheral_mscbus;

// DP6_26 input mux peripheral bus
input        [4:0] DP6_26_in_mux_peripheral_mscbus;

// DP6_27 input mux peripheral bus
input        [2:0] DP6_27_in_mux_peripheral_mscbus;

// DP7_0 input mux peripheral bus
input        [5:0] DP7_0_in_mux_peripheral_mscbus;

// DP7_1 input mux peripheral bus
input        [3:0] DP7_1_in_mux_peripheral_mscbus;

// DP7_1 output demux peripheral bus
output       [1:0] DP7_1_out_demux_peripheral_mscbus;

// DP7_2 input mux peripheral bus
input        [5:0] DP7_2_in_mux_peripheral_mscbus;

// DP7_3 input mux peripheral bus
input        [5:0] DP7_3_in_mux_peripheral_mscbus;

// DP7_4 input mux peripheral bus
input        [5:0] DP7_4_in_mux_peripheral_mscbus;

// DP7_5 input mux peripheral bus
input        [5:0] DP7_5_in_mux_peripheral_mscbus;

// DP7_6 input mux peripheral bus
input        [4:0] DP7_6_in_mux_peripheral_mscbus;

// DP7_6 output demux peripheral bus
output            DP7_6_out_demux_peripheral_mscbus;

// DP7_7 input mux peripheral bus
input        [4:0] DP7_7_in_mux_peripheral_mscbus;

// DP7_7 output demux peripheral bus
output       [1:0] DP7_7_out_demux_peripheral_mscbus;

// DP7_8 input mux peripheral bus
input        [5:0] DP7_8_in_mux_peripheral_mscbus;

// DP7_8 output demux peripheral bus
output            DP7_8_out_demux_peripheral_mscbus;

// DP7_9 input mux peripheral bus
input        [4:0] DP7_9_in_mux_peripheral_mscbus;

// DP7_9 output demux peripheral bus
output            DP7_9_out_demux_peripheral_mscbus;

// DP7_10 input mux peripheral bus
input             DP7_10_in_mux_peripheral_mscbus;

// DP7_10 output demux peripheral bus
output       [2:0] DP7_10_out_demux_peripheral_mscbus;

// DP7_11 input mux peripheral bus
input        [2:0] DP7_11_in_mux_peripheral_mscbus;

// DP7_11 output demux peripheral bus
output            DP7_11_out_demux_peripheral_mscbus;

// DP7_12 input mux peripheral bus
input        [1:0] DP7_12_in_mux_peripheral_mscbus;

// DP7_12 output demux peripheral bus
output       [1:0] DP7_12_out_demux_peripheral_mscbus;

// DP7_13 input mux peripheral bus
input        [1:0] DP7_13_in_mux_peripheral_mscbus;

// DP7_13 output demux peripheral bus
output       [1:0] DP7_13_out_demux_peripheral_mscbus;

// DP7_14 input mux peripheral bus
input             DP7_14_in_mux_peripheral_mscbus;

// DP7_14 output demux peripheral bus
output       [2:0] DP7_14_out_demux_peripheral_mscbus;

// DP7_15 input mux peripheral bus
input             DP7_15_in_mux_peripheral_mscbus;

// DP7_15 output demux peripheral bus
output       [1:0] DP7_15_out_demux_peripheral_mscbus;

// MP0_0 input mux peripheral bus
input        [2:0] MP0_0_in_mux_peripheral_mscbus;

// MP0_0 output demux peripheral bus
output            MP0_0_out_demux_peripheral_mscbus;

// MP0_1 input mux peripheral bus
input        [1:0] MP0_1_in_mux_peripheral_mscbus;

// MP0_1 output demux peripheral bus
output       [1:0] MP0_1_out_demux_peripheral_mscbus;

// MP0_2 input mux peripheral bus
input        [2:0] MP0_2_in_mux_peripheral_mscbus;

// MP0_2 output demux peripheral bus
output            MP0_2_out_demux_peripheral_mscbus;

// MP0_3 input mux peripheral bus
input        [1:0] MP0_3_in_mux_peripheral_mscbus;

// MP0_3 output demux peripheral bus
output       [1:0] MP0_3_out_demux_peripheral_mscbus;

// MP0_4 input mux peripheral bus
input        [2:0] MP0_4_in_mux_peripheral_mscbus;

// MP0_4 output demux peripheral bus
output            MP0_4_out_demux_peripheral_mscbus;

// MP0_5 output demux peripheral bus
output       [1:0] MP0_5_out_demux_peripheral_mscbus;

// MP0_6 input mux peripheral bus
input        [2:0] MP0_6_in_mux_peripheral_mscbus;

// MP0_6 output demux peripheral bus
output            MP0_6_out_demux_peripheral_mscbus;

// MP0_7 input mux peripheral bus
input        [1:0] MP0_7_in_mux_peripheral_mscbus;

// MP0_7 output demux peripheral bus
output       [1:0] MP0_7_out_demux_peripheral_mscbus;

// MP0_8 input mux peripheral bus
input        [3:0] MP0_8_in_mux_peripheral_mscbus;

// MP0_8 output demux peripheral bus
output            MP0_8_out_demux_peripheral_mscbus;

// MP0_9 input mux peripheral bus
input             MP0_9_in_mux_peripheral_mscbus;

// MP0_9 output demux peripheral bus
output       [2:0] MP0_9_out_demux_peripheral_mscbus;

// MP0_10 input mux peripheral bus
input        [2:0] MP0_10_in_mux_peripheral_mscbus;

// MP0_10 output demux peripheral bus
output            MP0_10_out_demux_peripheral_mscbus;

// MP0_11 output demux peripheral bus
output       [2:0] MP0_11_out_demux_peripheral_mscbus;

// MP0_12 input mux peripheral bus
input        [2:0] MP0_12_in_mux_peripheral_mscbus;

// MP0_12 output demux peripheral bus
output            MP0_12_out_demux_peripheral_mscbus;

// MP0_13 input mux peripheral bus
input             MP0_13_in_mux_peripheral_mscbus;

// MP0_13 output demux peripheral bus
output       [2:0] MP0_13_out_demux_peripheral_mscbus;

// MP0_14 input mux peripheral bus
input        [3:0] MP0_14_in_mux_peripheral_mscbus;

// MP0_15 input mux peripheral bus
input        [1:0] MP0_15_in_mux_peripheral_mscbus;

// MP0_15 output demux peripheral bus
output       [1:0] MP0_15_out_demux_peripheral_mscbus;

// MP0_16 input mux peripheral bus
input        [3:0] MP0_16_in_mux_peripheral_mscbus;

// MP0_17 output demux peripheral bus
output       [1:0] MP0_17_out_demux_peripheral_mscbus;

// MP0_18 input mux peripheral bus
input        [3:0] MP0_18_in_mux_peripheral_mscbus;

// MP0_19 input mux peripheral bus
input        [1:0] MP0_19_in_mux_peripheral_mscbus;

// MP0_19 output demux peripheral bus
output       [1:0] MP0_19_out_demux_peripheral_mscbus;

// MP0_20 input mux peripheral bus
input        [3:0] MP0_20_in_mux_peripheral_mscbus;

// MP0_21 input mux peripheral bus
input        [1:0] MP0_21_in_mux_peripheral_mscbus;

// MP0_21 output demux peripheral bus
output       [1:0] MP0_21_out_demux_peripheral_mscbus;

// MP0_22 input mux peripheral bus
input        [2:0] MP0_22_in_mux_peripheral_mscbus;

// MP0_23 input mux peripheral bus
input             MP0_23_in_mux_peripheral_mscbus;

// MP0_23 output demux peripheral bus
output            MP0_23_out_demux_peripheral_mscbus;

// MP0_24 input mux peripheral bus
input             MP0_24_in_mux_peripheral_mscbus;

// MP0_24 output demux peripheral bus
output       [1:0] MP0_24_out_demux_peripheral_mscbus;

// MP0_25 output demux peripheral bus
output       [2:0] MP0_25_out_demux_peripheral_mscbus;

// MP0_26 input mux peripheral bus
input        [1:0] MP0_26_in_mux_peripheral_mscbus;

// MP0_26 output demux peripheral bus
output            MP0_26_out_demux_peripheral_mscbus;

// MP0_27 output demux peripheral bus
output       [2:0] MP0_27_out_demux_peripheral_mscbus;

// MP0_28 input mux peripheral bus
input        [2:0] MP0_28_in_mux_peripheral_mscbus;

// MP0_29 output demux peripheral bus
output       [1:0] MP0_29_out_demux_peripheral_mscbus;

// MP0_30 input mux peripheral bus
input        [2:0] MP0_30_in_mux_peripheral_mscbus;

// MP0_31 input mux peripheral bus
input        [1:0] MP0_31_in_mux_peripheral_mscbus;

// MP0_31 output demux peripheral bus
output            MP0_31_out_demux_peripheral_mscbus;

// MP1_0 input mux peripheral bus
input        [2:0] MP1_0_in_mux_peripheral_mscbus;

// MP1_1 input mux peripheral bus
input        [1:0] MP1_1_in_mux_peripheral_mscbus;

// MP1_1 output demux peripheral bus
output            MP1_1_out_demux_peripheral_mscbus;

// MP1_2 input mux peripheral bus
input        [1:0] MP1_2_in_mux_peripheral_mscbus;

// MP1_2 output demux peripheral bus
output            MP1_2_out_demux_peripheral_mscbus;

// MP1_3 output demux peripheral bus
output       [1:0] MP1_3_out_demux_peripheral_mscbus;

// MP1_4 input mux peripheral bus
input             MP1_4_in_mux_peripheral_mscbus;

// MP1_4 output demux peripheral bus
output            MP1_4_out_demux_peripheral_mscbus;

// MP1_5 input mux peripheral bus
input             MP1_5_in_mux_peripheral_mscbus;

// MP1_5 output demux peripheral bus
output            MP1_5_out_demux_peripheral_mscbus;

// MP1_6 input mux peripheral bus
input             MP1_6_in_mux_peripheral_mscbus;

// MP1_6 output demux peripheral bus
output            MP1_6_out_demux_peripheral_mscbus;

// MP1_7 input mux peripheral bus
input             MP1_7_in_mux_peripheral_mscbus;

// MP1_7 output demux peripheral bus
output            MP1_7_out_demux_peripheral_mscbus;

// MP1_8 input mux peripheral bus
input             MP1_8_in_mux_peripheral_mscbus;

// MP1_8 output demux peripheral bus
output            MP1_8_out_demux_peripheral_mscbus;

// MP1_9 input mux peripheral bus
input             MP1_9_in_mux_peripheral_mscbus;

// MP1_9 output demux peripheral bus
output            MP1_9_out_demux_peripheral_mscbus;

// MP1_10 input mux peripheral bus
input        [1:0] MP1_10_in_mux_peripheral_mscbus;

// MP1_11 input mux peripheral bus
input        [1:0] MP1_11_in_mux_peripheral_mscbus;

// MP1_12 input mux peripheral bus
input             MP1_12_in_mux_peripheral_mscbus;

// MP1_13 input mux peripheral bus
input             MP1_13_in_mux_peripheral_mscbus;

// MP1_14 input mux peripheral bus
input             MP1_14_in_mux_peripheral_mscbus;

// MP1_15 input mux peripheral bus
input             MP1_15_in_mux_peripheral_mscbus;

// MP2_0 input mux peripheral bus
input        [2:0] MP2_0_in_mux_peripheral_mscbus;

// MP2_0 output demux peripheral bus
output            MP2_0_out_demux_peripheral_mscbus;

// MP2_1 input mux peripheral bus
input             MP2_1_in_mux_peripheral_mscbus;

// MP2_1 output demux peripheral bus
output       [2:0] MP2_1_out_demux_peripheral_mscbus;

// MP2_2 input mux peripheral bus
input        [2:0] MP2_2_in_mux_peripheral_mscbus;

// MP2_2 output demux peripheral bus
output            MP2_2_out_demux_peripheral_mscbus;

// MP2_3 input mux peripheral bus
input        [1:0] MP2_3_in_mux_peripheral_mscbus;

// MP2_3 output demux peripheral bus
output       [1:0] MP2_3_out_demux_peripheral_mscbus;

// MP2_4 input mux peripheral bus
input        [2:0] MP2_4_in_mux_peripheral_mscbus;

// MP2_4 output demux peripheral bus
output            MP2_4_out_demux_peripheral_mscbus;

// MP2_5 input mux peripheral bus
input        [1:0] MP2_5_in_mux_peripheral_mscbus;

// MP2_5 output demux peripheral bus
output       [1:0] MP2_5_out_demux_peripheral_mscbus;

// MP2_6 input mux peripheral bus
input        [2:0] MP2_6_in_mux_peripheral_mscbus;

// MP2_6 output demux peripheral bus
output            MP2_6_out_demux_peripheral_mscbus;

// MP2_7 input mux peripheral bus
input        [1:0] MP2_7_in_mux_peripheral_mscbus;

// MP2_7 output demux peripheral bus
output       [1:0] MP2_7_out_demux_peripheral_mscbus;

// MP2_8 input mux peripheral bus
input        [1:0] MP2_8_in_mux_peripheral_mscbus;

// MP2_8 output demux peripheral bus
output            MP2_8_out_demux_peripheral_mscbus;

// MP2_9 input mux peripheral bus
input             MP2_9_in_mux_peripheral_mscbus;

// MP2_9 output demux peripheral bus
output       [2:0] MP2_9_out_demux_peripheral_mscbus;

// MP2_10 input mux peripheral bus
input        [2:0] MP2_10_in_mux_peripheral_mscbus;

// MP2_10 output demux peripheral bus
output            MP2_10_out_demux_peripheral_mscbus;

// MP2_11 input mux peripheral bus
input        [1:0] MP2_11_in_mux_peripheral_mscbus;

// MP2_11 output demux peripheral bus
output       [1:0] MP2_11_out_demux_peripheral_mscbus;

// MP2_12 input mux peripheral bus
input        [1:0] MP2_12_in_mux_peripheral_mscbus;

// MP2_12 output demux peripheral bus
output       [1:0] MP2_12_out_demux_peripheral_mscbus;

// MP2_13 input mux peripheral bus
input             MP2_13_in_mux_peripheral_mscbus;

// MP2_13 output demux peripheral bus
output       [2:0] MP2_13_out_demux_peripheral_mscbus;

// MP2_14 input mux peripheral bus
input        [2:0] MP2_14_in_mux_peripheral_mscbus;

// MP2_14 output demux peripheral bus
output            MP2_14_out_demux_peripheral_mscbus;

// MP2_15 input mux peripheral bus
input             MP2_15_in_mux_peripheral_mscbus;

// MP2_15 output demux peripheral bus
output       [2:0] MP2_15_out_demux_peripheral_mscbus;

//======================================
// Signal Declarations
//======================================
wire      [6:0] DP0_0_in_mux_peripheral_mscbus;
wire      [4:0] DP0_10_in_mux_peripheral_mscbus;
wire      [4:0] DP0_11_in_mux_peripheral_mscbus;
wire      [4:0] DP0_12_in_mux_peripheral_mscbus;
wire      [4:0] DP0_13_in_mux_peripheral_mscbus;
wire            DP0_13_out_demux_peripheral_mscbus;
wire      [5:0] DP0_14_in_mux_peripheral_mscbus;
wire            DP0_14_out_demux_peripheral_mscbus;
wire      [5:0] DP0_15_in_mux_peripheral_mscbus;
wire            DP0_15_out_demux_peripheral_mscbus;
wire      [3:0] DP0_16_in_mux_peripheral_mscbus;
wire      [1:0] DP0_16_out_demux_peripheral_mscbus;
wire      [4:0] DP0_17_in_mux_peripheral_mscbus;
wire            DP0_17_out_demux_peripheral_mscbus;
wire      [4:0] DP0_18_in_mux_peripheral_mscbus;
wire            DP0_18_out_demux_peripheral_mscbus;
wire      [5:0] DP0_19_in_mux_peripheral_mscbus;
wire      [3:0] DP0_1_in_mux_peripheral_mscbus;
wire      [1:0] DP0_1_out_demux_peripheral_mscbus;
wire      [5:0] DP0_20_in_mux_peripheral_mscbus;
wire      [4:0] DP0_21_in_mux_peripheral_mscbus;
wire            DP0_21_out_demux_peripheral_mscbus;
wire      [3:0] DP0_22_in_mux_peripheral_mscbus;
wire      [1:0] DP0_22_out_demux_peripheral_mscbus;
wire      [3:0] DP0_23_in_mux_peripheral_mscbus;
wire      [1:0] DP0_23_out_demux_peripheral_mscbus;
wire      [3:0] DP0_24_in_mux_peripheral_mscbus;
wire      [1:0] DP0_24_out_demux_peripheral_mscbus;
wire      [4:0] DP0_25_in_mux_peripheral_mscbus;
wire            DP0_25_out_demux_peripheral_mscbus;
wire      [4:0] DP0_26_in_mux_peripheral_mscbus;
wire            DP0_26_out_demux_peripheral_mscbus;
wire      [4:0] DP0_27_in_mux_peripheral_mscbus;
wire            DP0_27_out_demux_peripheral_mscbus;
wire      [3:0] DP0_28_in_mux_peripheral_mscbus;
wire            DP0_28_out_demux_peripheral_mscbus;
wire      [2:0] DP0_29_in_mux_peripheral_mscbus;
wire      [1:0] DP0_29_out_demux_peripheral_mscbus;
wire      [5:0] DP0_2_in_mux_peripheral_mscbus;
wire      [2:0] DP0_30_in_mux_peripheral_mscbus;
wire      [1:0] DP0_30_out_demux_peripheral_mscbus;
wire      [3:0] DP0_31_in_mux_peripheral_mscbus;
wire            DP0_31_out_demux_peripheral_mscbus;
wire      [4:0] DP0_3_in_mux_peripheral_mscbus;
wire            DP0_3_out_demux_peripheral_mscbus;
wire      [5:0] DP0_4_in_mux_peripheral_mscbus;
wire      [4:0] DP0_5_in_mux_peripheral_mscbus;
wire            DP0_5_out_demux_peripheral_mscbus;
wire      [5:0] DP0_6_in_mux_peripheral_mscbus;
wire      [4:0] DP0_7_in_mux_peripheral_mscbus;
wire            DP0_7_out_demux_peripheral_mscbus;
wire      [4:0] DP0_8_in_mux_peripheral_mscbus;
wire            DP0_8_out_demux_peripheral_mscbus;
wire      [4:0] DP0_9_in_mux_peripheral_mscbus;
wire            DP0_9_out_demux_peripheral_mscbus;
wire      [2:0] DP1_0_in_mux_peripheral_mscbus;
wire      [1:0] DP1_0_out_demux_peripheral_mscbus;
wire      [1:0] DP1_10_in_mux_peripheral_mscbus;
wire      [1:0] DP1_10_out_demux_peripheral_mscbus;
wire      [1:0] DP1_11_in_mux_peripheral_mscbus;
wire      [1:0] DP1_11_out_demux_peripheral_mscbus;
wire      [1:0] DP1_12_in_mux_peripheral_mscbus;
wire            DP1_12_out_demux_peripheral_mscbus;
wire      [3:0] DP1_13_in_mux_peripheral_mscbus;
wire            DP1_13_out_demux_peripheral_mscbus;
wire      [1:0] DP1_14_in_mux_peripheral_mscbus;
wire      [2:0] DP1_14_out_demux_peripheral_mscbus;
wire      [3:0] DP1_15_in_mux_peripheral_mscbus;
wire            DP1_15_out_demux_peripheral_mscbus;
wire      [2:0] DP1_16_in_mux_peripheral_mscbus;
wire      [1:0] DP1_16_out_demux_peripheral_mscbus;
wire      [2:0] DP1_17_in_mux_peripheral_mscbus;
wire      [1:0] DP1_17_out_demux_peripheral_mscbus;
wire      [2:0] DP1_18_in_mux_peripheral_mscbus;
wire      [1:0] DP1_18_out_demux_peripheral_mscbus;
wire      [3:0] DP1_19_in_mux_peripheral_mscbus;
wire            DP1_19_out_demux_peripheral_mscbus;
wire      [2:0] DP1_1_in_mux_peripheral_mscbus;
wire      [1:0] DP1_1_out_demux_peripheral_mscbus;
wire      [2:0] DP1_20_in_mux_peripheral_mscbus;
wire      [1:0] DP1_20_out_demux_peripheral_mscbus;
wire      [3:0] DP1_21_in_mux_peripheral_mscbus;
wire            DP1_21_out_demux_peripheral_mscbus;
wire      [3:0] DP1_22_in_mux_peripheral_mscbus;
wire            DP1_22_out_demux_peripheral_mscbus;
wire      [2:0] DP1_23_in_mux_peripheral_mscbus;
wire            DP1_23_out_demux_peripheral_mscbus;
wire      [2:0] DP1_24_in_mux_peripheral_mscbus;
wire            DP1_24_out_demux_peripheral_mscbus;
wire      [4:0] DP1_25_in_mux_peripheral_mscbus;
wire      [4:0] DP1_26_in_mux_peripheral_mscbus;
wire      [4:0] DP1_27_in_mux_peripheral_mscbus;
wire      [3:0] DP1_28_in_mux_peripheral_mscbus;
wire            DP1_28_out_demux_peripheral_mscbus;
wire      [3:0] DP1_29_in_mux_peripheral_mscbus;
wire            DP1_29_out_demux_peripheral_mscbus;
wire      [2:0] DP1_2_in_mux_peripheral_mscbus;
wire      [1:0] DP1_2_out_demux_peripheral_mscbus;
wire      [3:0] DP1_30_in_mux_peripheral_mscbus;
wire            DP1_30_out_demux_peripheral_mscbus;
wire      [2:0] DP1_31_in_mux_peripheral_mscbus;
wire      [1:0] DP1_31_out_demux_peripheral_mscbus;
wire      [3:0] DP1_3_in_mux_peripheral_mscbus;
wire            DP1_3_out_demux_peripheral_mscbus;
wire      [3:0] DP1_4_in_mux_peripheral_mscbus;
wire            DP1_4_out_demux_peripheral_mscbus;
wire      [3:0] DP1_5_in_mux_peripheral_mscbus;
wire            DP1_5_out_demux_peripheral_mscbus;
wire      [2:0] DP1_6_in_mux_peripheral_mscbus;
wire      [1:0] DP1_6_out_demux_peripheral_mscbus;
wire      [3:0] DP1_7_in_mux_peripheral_mscbus;
wire            DP1_7_out_demux_peripheral_mscbus;
wire      [2:0] DP1_8_in_mux_peripheral_mscbus;
wire            DP1_8_out_demux_peripheral_mscbus;
wire      [2:0] DP1_9_in_mux_peripheral_mscbus;
wire            DP1_9_out_demux_peripheral_mscbus;
wire      [3:0] DP2_0_in_mux_peripheral_mscbus;
wire            DP2_0_out_demux_peripheral_mscbus;
wire      [3:0] DP2_10_in_mux_peripheral_mscbus;
wire      [2:0] DP2_11_in_mux_peripheral_mscbus;
wire      [3:0] DP2_12_in_mux_peripheral_mscbus;
wire            DP2_12_out_demux_peripheral_mscbus;
wire      [2:0] DP2_13_in_mux_peripheral_mscbus;
wire            DP2_13_out_demux_peripheral_mscbus;
wire      [3:0] DP2_14_in_mux_peripheral_mscbus;
wire      [2:0] DP2_15_in_mux_peripheral_mscbus;
wire            DP2_15_out_demux_peripheral_mscbus;
wire      [2:0] DP2_16_in_mux_peripheral_mscbus;
wire            DP2_16_out_demux_peripheral_mscbus;
wire      [2:0] DP2_17_in_mux_peripheral_mscbus;
wire            DP2_17_out_demux_peripheral_mscbus;
wire      [3:0] DP2_18_in_mux_peripheral_mscbus;
wire      [3:0] DP2_19_in_mux_peripheral_mscbus;
wire      [3:0] DP2_1_in_mux_peripheral_mscbus;
wire      [2:0] DP2_20_in_mux_peripheral_mscbus;
wire            DP2_20_out_demux_peripheral_mscbus;
wire      [5:0] DP2_21_in_mux_peripheral_mscbus;
wire      [4:0] DP2_22_in_mux_peripheral_mscbus;
wire            DP2_22_out_demux_peripheral_mscbus;
wire      [5:0] DP2_23_in_mux_peripheral_mscbus;
wire            DP2_23_out_demux_peripheral_mscbus;
wire      [4:0] DP2_24_in_mux_peripheral_mscbus;
wire      [1:0] DP2_24_out_demux_peripheral_mscbus;
wire      [5:0] DP2_25_in_mux_peripheral_mscbus;
wire      [3:0] DP2_26_in_mux_peripheral_mscbus;
wire      [1:0] DP2_26_out_demux_peripheral_mscbus;
wire      [4:0] DP2_27_in_mux_peripheral_mscbus;
wire            DP2_27_out_demux_peripheral_mscbus;
wire      [2:0] DP2_28_in_mux_peripheral_mscbus;
wire      [2:0] DP2_28_out_demux_peripheral_mscbus;
wire      [4:0] DP2_29_in_mux_peripheral_mscbus;
wire            DP2_29_out_demux_peripheral_mscbus;
wire      [3:0] DP2_2_in_mux_peripheral_mscbus;
wire            DP2_2_out_demux_peripheral_mscbus;
wire      [3:0] DP2_30_in_mux_peripheral_mscbus;
wire      [1:0] DP2_30_out_demux_peripheral_mscbus;
wire      [4:0] DP2_31_in_mux_peripheral_mscbus;
wire            DP2_31_out_demux_peripheral_mscbus;
wire      [3:0] DP2_3_in_mux_peripheral_mscbus;
wire            DP2_3_out_demux_peripheral_mscbus;
wire      [3:0] DP2_4_in_mux_peripheral_mscbus;
wire      [3:0] DP2_5_in_mux_peripheral_mscbus;
wire      [2:0] DP2_6_in_mux_peripheral_mscbus;
wire            DP2_6_out_demux_peripheral_mscbus;
wire      [3:0] DP2_7_in_mux_peripheral_mscbus;
wire      [3:0] DP2_8_in_mux_peripheral_mscbus;
wire      [3:0] DP2_9_in_mux_peripheral_mscbus;
wire      [3:0] DP3_0_in_mux_peripheral_mscbus;
wire      [1:0] DP3_0_out_demux_peripheral_mscbus;
wire      [2:0] DP3_10_in_mux_peripheral_mscbus;
wire      [2:0] DP3_10_out_demux_peripheral_mscbus;
wire      [3:0] DP3_11_in_mux_peripheral_mscbus;
wire      [1:0] DP3_11_out_demux_peripheral_mscbus;
wire      [5:0] DP3_12_in_mux_peripheral_mscbus;
wire      [3:0] DP3_13_in_mux_peripheral_mscbus;
wire      [1:0] DP3_13_out_demux_peripheral_mscbus;
wire      [5:0] DP3_14_in_mux_peripheral_mscbus;
wire      [4:0] DP3_15_in_mux_peripheral_mscbus;
wire            DP3_15_out_demux_peripheral_mscbus;
wire      [4:0] DP3_16_in_mux_peripheral_mscbus;
wire            DP3_16_out_demux_peripheral_mscbus;
wire      [3:0] DP3_17_in_mux_peripheral_mscbus;
wire      [1:0] DP3_17_out_demux_peripheral_mscbus;
wire      [5:0] DP3_18_in_mux_peripheral_mscbus;
wire      [5:0] DP3_19_in_mux_peripheral_mscbus;
wire      [3:0] DP3_1_in_mux_peripheral_mscbus;
wire      [1:0] DP3_1_out_demux_peripheral_mscbus;
wire      [5:0] DP3_20_in_mux_peripheral_mscbus;
wire      [6:0] DP3_21_in_mux_peripheral_mscbus;
wire      [6:0] DP3_22_in_mux_peripheral_mscbus;
wire      [6:0] DP3_23_in_mux_peripheral_mscbus;
wire      [4:0] DP3_24_in_mux_peripheral_mscbus;
wire      [1:0] DP3_24_out_demux_peripheral_mscbus;
wire      [5:0] DP3_25_in_mux_peripheral_mscbus;
wire            DP3_25_out_demux_peripheral_mscbus;
wire      [4:0] DP3_26_in_mux_peripheral_mscbus;
wire      [1:0] DP3_26_out_demux_peripheral_mscbus;
wire      [4:0] DP3_27_in_mux_peripheral_mscbus;
wire      [1:0] DP3_27_out_demux_peripheral_mscbus;
wire      [4:0] DP3_28_in_mux_peripheral_mscbus;
wire      [1:0] DP3_28_out_demux_peripheral_mscbus;
wire      [4:0] DP3_29_in_mux_peripheral_mscbus;
wire      [4:0] DP3_2_in_mux_peripheral_mscbus;
wire            DP3_2_out_demux_peripheral_mscbus;
wire      [4:0] DP3_30_in_mux_peripheral_mscbus;
wire            DP3_30_out_demux_peripheral_mscbus;
wire      [2:0] DP3_31_in_mux_peripheral_mscbus;
wire      [2:0] DP3_31_out_demux_peripheral_mscbus;
wire      [2:0] DP3_3_in_mux_peripheral_mscbus;
wire      [2:0] DP3_3_out_demux_peripheral_mscbus;
wire      [4:0] DP3_4_in_mux_peripheral_mscbus;
wire            DP3_4_out_demux_peripheral_mscbus;
wire      [3:0] DP3_5_in_mux_peripheral_mscbus;
wire            DP3_5_out_demux_peripheral_mscbus;
wire      [3:0] DP3_6_in_mux_peripheral_mscbus;
wire            DP3_6_out_demux_peripheral_mscbus;
wire      [3:0] DP3_7_in_mux_peripheral_mscbus;
wire            DP3_7_out_demux_peripheral_mscbus;
wire      [4:0] DP3_8_in_mux_peripheral_mscbus;
wire            DP3_8_out_demux_peripheral_mscbus;
wire      [3:0] DP3_9_in_mux_peripheral_mscbus;
wire      [1:0] DP3_9_out_demux_peripheral_mscbus;
wire      [3:0] DP4_0_in_mux_peripheral_mscbus;
wire            DP4_0_out_demux_peripheral_mscbus;
wire      [4:0] DP4_10_in_mux_peripheral_mscbus;
wire      [1:0] DP4_10_out_demux_peripheral_mscbus;
wire      [5:0] DP4_11_in_mux_peripheral_mscbus;
wire            DP4_11_out_demux_peripheral_mscbus;
wire      [4:0] DP4_12_in_mux_peripheral_mscbus;
wire      [1:0] DP4_12_out_demux_peripheral_mscbus;
wire      [4:0] DP4_13_in_mux_peripheral_mscbus;
wire      [1:0] DP4_13_out_demux_peripheral_mscbus;
wire      [3:0] DP4_14_in_mux_peripheral_mscbus;
wire            DP4_14_out_demux_peripheral_mscbus;
wire      [3:0] DP4_15_in_mux_peripheral_mscbus;
wire      [2:0] DP4_15_out_demux_peripheral_mscbus;
wire      [3:0] DP4_16_in_mux_peripheral_mscbus;
wire      [2:0] DP4_16_out_demux_peripheral_mscbus;
wire      [3:0] DP4_17_in_mux_peripheral_mscbus;
wire      [2:0] DP4_17_out_demux_peripheral_mscbus;
wire      [1:0] DP4_18_in_mux_peripheral_mscbus;
wire      [1:0] DP4_18_out_demux_peripheral_mscbus;
wire      [2:0] DP4_19_in_mux_peripheral_mscbus;
wire      [2:0] DP4_1_in_mux_peripheral_mscbus;
wire      [1:0] DP4_1_out_demux_peripheral_mscbus;
wire      [5:0] DP4_20_in_mux_peripheral_mscbus;
wire      [5:0] DP4_21_in_mux_peripheral_mscbus;
wire      [4:0] DP4_22_in_mux_peripheral_mscbus;
wire            DP4_22_out_demux_peripheral_mscbus;
wire      [4:0] DP4_23_in_mux_peripheral_mscbus;
wire      [4:0] DP4_24_in_mux_peripheral_mscbus;
wire      [2:0] DP4_25_in_mux_peripheral_mscbus;
wire            DP4_25_out_demux_peripheral_mscbus;
wire      [3:0] DP4_26_in_mux_peripheral_mscbus;
wire      [3:0] DP4_27_in_mux_peripheral_mscbus;
wire            DP4_27_out_demux_peripheral_mscbus;
wire      [4:0] DP4_28_in_mux_peripheral_mscbus;
wire            DP4_28_out_demux_peripheral_mscbus;
wire      [2:0] DP4_29_in_mux_peripheral_mscbus;
wire      [1:0] DP4_29_out_demux_peripheral_mscbus;
wire      [3:0] DP4_2_in_mux_peripheral_mscbus;
wire            DP4_2_out_demux_peripheral_mscbus;
wire      [3:0] DP4_30_in_mux_peripheral_mscbus;
wire            DP4_30_out_demux_peripheral_mscbus;
wire      [2:0] DP4_31_in_mux_peripheral_mscbus;
wire      [1:0] DP4_31_out_demux_peripheral_mscbus;
wire      [3:0] DP4_3_in_mux_peripheral_mscbus;
wire            DP4_3_out_demux_peripheral_mscbus;
wire      [2:0] DP4_4_in_mux_peripheral_mscbus;
wire      [1:0] DP4_4_out_demux_peripheral_mscbus;
wire      [4:0] DP4_5_in_mux_peripheral_mscbus;
wire      [5:0] DP4_6_in_mux_peripheral_mscbus;
wire      [1:0] DP4_6_out_demux_peripheral_mscbus;
wire      [5:0] DP4_7_in_mux_peripheral_mscbus;
wire            DP4_7_out_demux_peripheral_mscbus;
wire      [6:0] DP4_8_in_mux_peripheral_mscbus;
wire      [4:0] DP4_9_in_mux_peripheral_mscbus;
wire      [1:0] DP4_9_out_demux_peripheral_mscbus;
wire      [6:0] DP5_0_in_mux_peripheral_mscbus;
wire      [4:0] DP5_10_in_mux_peripheral_mscbus;
wire      [1:0] DP5_10_out_demux_peripheral_mscbus;
wire      [3:0] DP5_11_in_mux_peripheral_mscbus;
wire      [2:0] DP5_11_out_demux_peripheral_mscbus;
wire      [4:0] DP5_12_in_mux_peripheral_mscbus;
wire      [1:0] DP5_12_out_demux_peripheral_mscbus;
wire      [4:0] DP5_13_in_mux_peripheral_mscbus;
wire      [1:0] DP5_13_out_demux_peripheral_mscbus;
wire      [5:0] DP5_14_in_mux_peripheral_mscbus;
wire      [4:0] DP5_15_in_mux_peripheral_mscbus;
wire            DP5_15_out_demux_peripheral_mscbus;
wire      [4:0] DP5_16_in_mux_peripheral_mscbus;
wire            DP5_16_out_demux_peripheral_mscbus;
wire      [4:0] DP5_17_in_mux_peripheral_mscbus;
wire            DP5_17_out_demux_peripheral_mscbus;
wire      [4:0] DP5_18_in_mux_peripheral_mscbus;
wire      [3:0] DP5_19_in_mux_peripheral_mscbus;
wire            DP5_19_out_demux_peripheral_mscbus;
wire      [4:0] DP5_1_in_mux_peripheral_mscbus;
wire            DP5_1_out_demux_peripheral_mscbus;
wire      [5:0] DP5_20_in_mux_peripheral_mscbus;
wire      [4:0] DP5_21_in_mux_peripheral_mscbus;
wire            DP5_21_out_demux_peripheral_mscbus;
wire      [3:0] DP5_22_in_mux_peripheral_mscbus;
wire      [1:0] DP5_22_out_demux_peripheral_mscbus;
wire      [4:0] DP5_23_in_mux_peripheral_mscbus;
wire            DP5_23_out_demux_peripheral_mscbus;
wire      [4:0] DP5_24_in_mux_peripheral_mscbus;
wire            DP5_24_out_demux_peripheral_mscbus;
wire      [3:0] DP5_25_in_mux_peripheral_mscbus;
wire            DP5_25_out_demux_peripheral_mscbus;
wire      [5:0] DP5_26_in_mux_peripheral_mscbus;
wire            DP5_26_out_demux_peripheral_mscbus;
wire      [7:0] DP5_27_in_mux_peripheral_mscbus;
wire      [5:0] DP5_28_in_mux_peripheral_mscbus;
wire      [1:0] DP5_28_out_demux_peripheral_mscbus;
wire      [6:0] DP5_29_in_mux_peripheral_mscbus;
wire            DP5_29_out_demux_peripheral_mscbus;
wire      [4:0] DP5_2_in_mux_peripheral_mscbus;
wire            DP5_2_out_demux_peripheral_mscbus;
wire      [4:0] DP5_30_in_mux_peripheral_mscbus;
wire      [2:0] DP5_30_out_demux_peripheral_mscbus;
wire      [6:0] DP5_31_in_mux_peripheral_mscbus;
wire            DP5_31_out_demux_peripheral_mscbus;
wire      [4:0] DP5_3_in_mux_peripheral_mscbus;
wire            DP5_3_out_demux_peripheral_mscbus;
wire      [4:0] DP5_4_in_mux_peripheral_mscbus;
wire      [1:0] DP5_4_out_demux_peripheral_mscbus;
wire      [4:0] DP5_5_in_mux_peripheral_mscbus;
wire      [1:0] DP5_5_out_demux_peripheral_mscbus;
wire      [6:0] DP5_6_in_mux_peripheral_mscbus;
wire            DP5_6_out_demux_peripheral_mscbus;
wire      [6:0] DP5_7_in_mux_peripheral_mscbus;
wire      [5:0] DP5_8_in_mux_peripheral_mscbus;
wire            DP5_8_out_demux_peripheral_mscbus;
wire      [2:0] DP5_9_in_mux_peripheral_mscbus;
wire      [3:0] DP5_9_out_demux_peripheral_mscbus;
wire      [4:0] DP6_0_in_mux_peripheral_mscbus;
wire      [2:0] DP6_0_out_demux_peripheral_mscbus;
wire      [4:0] DP6_10_in_mux_peripheral_mscbus;
wire            DP6_10_out_demux_peripheral_mscbus;
wire      [5:0] DP6_11_in_mux_peripheral_mscbus;
wire      [5:0] DP6_12_in_mux_peripheral_mscbus;
wire            DP6_12_out_demux_peripheral_mscbus;
wire      [5:0] DP6_13_in_mux_peripheral_mscbus;
wire      [1:0] DP6_13_out_demux_peripheral_mscbus;
wire      [5:0] DP6_14_in_mux_peripheral_mscbus;
wire            DP6_14_out_demux_peripheral_mscbus;
wire      [4:0] DP6_15_in_mux_peripheral_mscbus;
wire      [1:0] DP6_15_out_demux_peripheral_mscbus;
wire      [5:0] DP6_16_in_mux_peripheral_mscbus;
wire            DP6_16_out_demux_peripheral_mscbus;
wire      [6:0] DP6_17_in_mux_peripheral_mscbus;
wire      [6:0] DP6_18_in_mux_peripheral_mscbus;
wire            DP6_18_out_demux_peripheral_mscbus;
wire      [4:0] DP6_19_in_mux_peripheral_mscbus;
wire      [1:0] DP6_19_out_demux_peripheral_mscbus;
wire      [4:0] DP6_1_in_mux_peripheral_mscbus;
wire      [1:0] DP6_1_out_demux_peripheral_mscbus;
wire      [6:0] DP6_20_in_mux_peripheral_mscbus;
wire      [3:0] DP6_21_in_mux_peripheral_mscbus;
wire      [2:0] DP6_21_out_demux_peripheral_mscbus;
wire      [4:0] DP6_22_in_mux_peripheral_mscbus;
wire      [1:0] DP6_22_out_demux_peripheral_mscbus;
wire      [5:0] DP6_23_in_mux_peripheral_mscbus;
wire            DP6_23_out_demux_peripheral_mscbus;
wire      [5:0] DP6_24_in_mux_peripheral_mscbus;
wire            DP6_24_out_demux_peripheral_mscbus;
wire      [4:0] DP6_25_in_mux_peripheral_mscbus;
wire      [1:0] DP6_25_out_demux_peripheral_mscbus;
wire      [4:0] DP6_26_in_mux_peripheral_mscbus;
wire      [2:0] DP6_27_in_mux_peripheral_mscbus;
wire      [4:0] DP6_2_in_mux_peripheral_mscbus;
wire      [2:0] DP6_2_out_demux_peripheral_mscbus;
wire      [6:0] DP6_3_in_mux_peripheral_mscbus;
wire            DP6_3_out_demux_peripheral_mscbus;
wire      [4:0] DP6_4_in_mux_peripheral_mscbus;
wire      [1:0] DP6_4_out_demux_peripheral_mscbus;
wire      [4:0] DP6_5_in_mux_peripheral_mscbus;
wire      [1:0] DP6_5_out_demux_peripheral_mscbus;
wire      [5:0] DP6_6_in_mux_peripheral_mscbus;
wire            DP6_6_out_demux_peripheral_mscbus;
wire      [5:0] DP6_7_in_mux_peripheral_mscbus;
wire            DP6_7_out_demux_peripheral_mscbus;
wire      [3:0] DP6_8_in_mux_peripheral_mscbus;
wire      [1:0] DP6_8_out_demux_peripheral_mscbus;
wire      [4:0] DP6_9_in_mux_peripheral_mscbus;
wire            DP6_9_out_demux_peripheral_mscbus;
wire      [5:0] DP7_0_in_mux_peripheral_mscbus;
wire            DP7_10_in_mux_peripheral_mscbus;
wire      [2:0] DP7_10_out_demux_peripheral_mscbus;
wire      [2:0] DP7_11_in_mux_peripheral_mscbus;
wire            DP7_11_out_demux_peripheral_mscbus;
wire      [1:0] DP7_12_in_mux_peripheral_mscbus;
wire      [1:0] DP7_12_out_demux_peripheral_mscbus;
wire      [1:0] DP7_13_in_mux_peripheral_mscbus;
wire      [1:0] DP7_13_out_demux_peripheral_mscbus;
wire            DP7_14_in_mux_peripheral_mscbus;
wire      [2:0] DP7_14_out_demux_peripheral_mscbus;
wire            DP7_15_in_mux_peripheral_mscbus;
wire      [1:0] DP7_15_out_demux_peripheral_mscbus;
wire      [3:0] DP7_1_in_mux_peripheral_mscbus;
wire      [1:0] DP7_1_out_demux_peripheral_mscbus;
wire      [5:0] DP7_2_in_mux_peripheral_mscbus;
wire      [5:0] DP7_3_in_mux_peripheral_mscbus;
wire      [5:0] DP7_4_in_mux_peripheral_mscbus;
wire      [5:0] DP7_5_in_mux_peripheral_mscbus;
wire      [4:0] DP7_6_in_mux_peripheral_mscbus;
wire            DP7_6_out_demux_peripheral_mscbus;
wire      [4:0] DP7_7_in_mux_peripheral_mscbus;
wire      [1:0] DP7_7_out_demux_peripheral_mscbus;
wire      [5:0] DP7_8_in_mux_peripheral_mscbus;
wire            DP7_8_out_demux_peripheral_mscbus;
wire      [4:0] DP7_9_in_mux_peripheral_mscbus;
wire            DP7_9_out_demux_peripheral_mscbus;
wire      [2:0] MP0_0_in_mux_peripheral_mscbus;
wire            MP0_0_out_demux_peripheral_mscbus;
wire      [2:0] MP0_10_in_mux_peripheral_mscbus;
wire            MP0_10_out_demux_peripheral_mscbus;
wire      [2:0] MP0_11_out_demux_peripheral_mscbus;
wire      [2:0] MP0_12_in_mux_peripheral_mscbus;
wire            MP0_12_out_demux_peripheral_mscbus;
wire            MP0_13_in_mux_peripheral_mscbus;
wire      [2:0] MP0_13_out_demux_peripheral_mscbus;
wire      [3:0] MP0_14_in_mux_peripheral_mscbus;
wire      [1:0] MP0_15_in_mux_peripheral_mscbus;
wire      [1:0] MP0_15_out_demux_peripheral_mscbus;
wire      [3:0] MP0_16_in_mux_peripheral_mscbus;
wire      [1:0] MP0_17_out_demux_peripheral_mscbus;
wire      [3:0] MP0_18_in_mux_peripheral_mscbus;
wire      [1:0] MP0_19_in_mux_peripheral_mscbus;
wire      [1:0] MP0_19_out_demux_peripheral_mscbus;
wire      [1:0] MP0_1_in_mux_peripheral_mscbus;
wire      [1:0] MP0_1_out_demux_peripheral_mscbus;
wire      [3:0] MP0_20_in_mux_peripheral_mscbus;
wire      [1:0] MP0_21_in_mux_peripheral_mscbus;
wire      [1:0] MP0_21_out_demux_peripheral_mscbus;
wire      [2:0] MP0_22_in_mux_peripheral_mscbus;
wire            MP0_23_in_mux_peripheral_mscbus;
wire            MP0_23_out_demux_peripheral_mscbus;
wire            MP0_24_in_mux_peripheral_mscbus;
wire      [1:0] MP0_24_out_demux_peripheral_mscbus;
wire      [2:0] MP0_25_out_demux_peripheral_mscbus;
wire      [1:0] MP0_26_in_mux_peripheral_mscbus;
wire            MP0_26_out_demux_peripheral_mscbus;
wire      [2:0] MP0_27_out_demux_peripheral_mscbus;
wire      [2:0] MP0_28_in_mux_peripheral_mscbus;
wire      [1:0] MP0_29_out_demux_peripheral_mscbus;
wire      [2:0] MP0_2_in_mux_peripheral_mscbus;
wire            MP0_2_out_demux_peripheral_mscbus;
wire      [2:0] MP0_30_in_mux_peripheral_mscbus;
wire      [1:0] MP0_31_in_mux_peripheral_mscbus;
wire            MP0_31_out_demux_peripheral_mscbus;
wire      [1:0] MP0_3_in_mux_peripheral_mscbus;
wire      [1:0] MP0_3_out_demux_peripheral_mscbus;
wire      [2:0] MP0_4_in_mux_peripheral_mscbus;
wire            MP0_4_out_demux_peripheral_mscbus;
wire      [1:0] MP0_5_out_demux_peripheral_mscbus;
wire      [2:0] MP0_6_in_mux_peripheral_mscbus;
wire            MP0_6_out_demux_peripheral_mscbus;
wire      [1:0] MP0_7_in_mux_peripheral_mscbus;
wire      [1:0] MP0_7_out_demux_peripheral_mscbus;
wire      [3:0] MP0_8_in_mux_peripheral_mscbus;
wire            MP0_8_out_demux_peripheral_mscbus;
wire            MP0_9_in_mux_peripheral_mscbus;
wire      [2:0] MP0_9_out_demux_peripheral_mscbus;
wire      [2:0] MP1_0_in_mux_peripheral_mscbus;
wire      [1:0] MP1_10_in_mux_peripheral_mscbus;
wire      [1:0] MP1_11_in_mux_peripheral_mscbus;
wire            MP1_12_in_mux_peripheral_mscbus;
wire            MP1_13_in_mux_peripheral_mscbus;
wire            MP1_14_in_mux_peripheral_mscbus;
wire            MP1_15_in_mux_peripheral_mscbus;
wire      [1:0] MP1_1_in_mux_peripheral_mscbus;
wire            MP1_1_out_demux_peripheral_mscbus;
wire      [1:0] MP1_2_in_mux_peripheral_mscbus;
wire            MP1_2_out_demux_peripheral_mscbus;
wire      [1:0] MP1_3_out_demux_peripheral_mscbus;
wire            MP1_4_in_mux_peripheral_mscbus;
wire            MP1_4_out_demux_peripheral_mscbus;
wire            MP1_5_in_mux_peripheral_mscbus;
wire            MP1_5_out_demux_peripheral_mscbus;
wire            MP1_6_in_mux_peripheral_mscbus;
wire            MP1_6_out_demux_peripheral_mscbus;
wire            MP1_7_in_mux_peripheral_mscbus;
wire            MP1_7_out_demux_peripheral_mscbus;
wire            MP1_8_in_mux_peripheral_mscbus;
wire            MP1_8_out_demux_peripheral_mscbus;
wire            MP1_9_in_mux_peripheral_mscbus;
wire            MP1_9_out_demux_peripheral_mscbus;
wire      [2:0] MP2_0_in_mux_peripheral_mscbus;
wire            MP2_0_out_demux_peripheral_mscbus;
wire      [2:0] MP2_10_in_mux_peripheral_mscbus;
wire            MP2_10_out_demux_peripheral_mscbus;
wire      [1:0] MP2_11_in_mux_peripheral_mscbus;
wire      [1:0] MP2_11_out_demux_peripheral_mscbus;
wire      [1:0] MP2_12_in_mux_peripheral_mscbus;
wire      [1:0] MP2_12_out_demux_peripheral_mscbus;
wire            MP2_13_in_mux_peripheral_mscbus;
wire      [2:0] MP2_13_out_demux_peripheral_mscbus;
wire      [2:0] MP2_14_in_mux_peripheral_mscbus;
wire            MP2_14_out_demux_peripheral_mscbus;
wire            MP2_15_in_mux_peripheral_mscbus;
wire      [2:0] MP2_15_out_demux_peripheral_mscbus;
wire            MP2_1_in_mux_peripheral_mscbus;
wire      [2:0] MP2_1_out_demux_peripheral_mscbus;
wire      [2:0] MP2_2_in_mux_peripheral_mscbus;
wire            MP2_2_out_demux_peripheral_mscbus;
wire      [1:0] MP2_3_in_mux_peripheral_mscbus;
wire      [1:0] MP2_3_out_demux_peripheral_mscbus;
wire      [2:0] MP2_4_in_mux_peripheral_mscbus;
wire            MP2_4_out_demux_peripheral_mscbus;
wire      [1:0] MP2_5_in_mux_peripheral_mscbus;
wire      [1:0] MP2_5_out_demux_peripheral_mscbus;
wire      [2:0] MP2_6_in_mux_peripheral_mscbus;
wire            MP2_6_out_demux_peripheral_mscbus;
wire      [1:0] MP2_7_in_mux_peripheral_mscbus;
wire      [1:0] MP2_7_out_demux_peripheral_mscbus;
wire      [1:0] MP2_8_in_mux_peripheral_mscbus;
wire            MP2_8_out_demux_peripheral_mscbus;
wire            MP2_9_in_mux_peripheral_mscbus;
wire      [2:0] MP2_9_out_demux_peripheral_mscbus;
wire     [31:0] ap_GP_DATA_IN_out_mscbus;
wire     [31:0] ap_amsel_out_mscbus;
wire     [31:0] ap_async_in_from_pad_mscbus;
wire     [31:0] ap_data_out_2_pinmux_mscbus;
wire     [31:0] ap_dir_out_mscbus;
wire     [31:0] ap_ds0_out_mscbus;
wire     [31:0] ap_ds1_out_mscbus;
wire     [31:0] ap_glitch_filter_bypass_out_mscbus;
wire     [63:0] ap_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] ap_gpio_out_2_buf_mscbus;
wire     [31:0] ap_gpio_out_en_2_buf_mscbus;
wire   [1023:0] ap_in_function_en_out_mscbus;
wire     [31:0] ap_in_termination_en_out_mscbus;
wire     [31:0] ap_inena_out_mscbus;
wire     [31:0] ap_lvds_en_ctrl_out_mscbus;
wire     [31:0] ap_mode0_out_mscbus;
wire     [31:0] ap_mode1_out_mscbus;
wire    [255:0] ap_pes_en_out_mscbus;
wire     [31:0] ap_pes_in_en_out_mscbus;
wire     [63:0] ap_pes_safeval_out_mscbus;
wire    [159:0] ap_pinmux_muxsel_out_mscbus;
wire     [31:0] ap_pinmuxdata_2_gpio_mscbus;
wire     [31:0] ap_pinmuxen_2_gpio_mscbus;
wire     [31:0] ap_pull_en_out_mscbus;
wire     [31:0] ap_pull_type_out_mscbus;
wire     [31:0] ap_schmitt_out_mscbus;
wire     [31:0] ap_slew_out_mscbus;
wire     [31:0] dp0_GP_DATA_IN_out_mscbus;
wire     [31:0] dp0_amsel_out_mscbus;
wire     [31:0] dp0_async_in_from_pad_mscbus;
wire     [31:0] dp0_data_out_2_pinmux_mscbus;
wire     [31:0] dp0_dir_out_mscbus;
wire     [31:0] dp0_ds0_out_mscbus;
wire     [31:0] dp0_ds1_out_mscbus;
wire     [31:0] dp0_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp0_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp0_gpio_out_2_buf_mscbus;
wire     [31:0] dp0_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp0_in_function_en_out_mscbus;
wire     [31:0] dp0_in_termination_en_out_mscbus;
wire     [31:0] dp0_inena_out_mscbus;
wire     [31:0] dp0_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp0_mode0_out_mscbus;
wire     [31:0] dp0_mode1_out_mscbus;
wire    [255:0] dp0_pes_en_out_mscbus;
wire     [31:0] dp0_pes_in_en_out_mscbus;
wire     [63:0] dp0_pes_safeval_out_mscbus;
wire    [159:0] dp0_pinmux_muxsel_out_mscbus;
wire     [31:0] dp0_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp0_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp0_pull_en_out_mscbus;
wire     [31:0] dp0_pull_type_out_mscbus;
wire     [31:0] dp0_schmitt_out_mscbus;
wire     [31:0] dp0_slew_out_mscbus;
wire     [31:0] dp1_GP_DATA_IN_out_mscbus;
wire     [31:0] dp1_amsel_out_mscbus;
wire     [31:0] dp1_async_in_from_pad_mscbus;
wire     [31:0] dp1_data_out_2_pinmux_mscbus;
wire     [31:0] dp1_dir_out_mscbus;
wire     [31:0] dp1_ds0_out_mscbus;
wire     [31:0] dp1_ds1_out_mscbus;
wire     [31:0] dp1_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp1_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp1_gpio_out_2_buf_mscbus;
wire     [31:0] dp1_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp1_in_function_en_out_mscbus;
wire     [31:0] dp1_in_termination_en_out_mscbus;
wire     [31:0] dp1_inena_out_mscbus;
wire     [31:0] dp1_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp1_mode0_out_mscbus;
wire     [31:0] dp1_mode1_out_mscbus;
wire    [255:0] dp1_pes_en_out_mscbus;
wire     [31:0] dp1_pes_in_en_out_mscbus;
wire     [63:0] dp1_pes_safeval_out_mscbus;
wire    [159:0] dp1_pinmux_muxsel_out_mscbus;
wire     [31:0] dp1_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp1_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp1_pull_en_out_mscbus;
wire     [31:0] dp1_pull_type_out_mscbus;
wire     [31:0] dp1_schmitt_out_mscbus;
wire     [31:0] dp1_slew_out_mscbus;
wire     [31:0] dp2_GP_DATA_IN_out_mscbus;
wire     [31:0] dp2_amsel_out_mscbus;
wire     [31:0] dp2_async_in_from_pad_mscbus;
wire     [31:0] dp2_data_out_2_pinmux_mscbus;
wire     [31:0] dp2_dir_out_mscbus;
wire     [31:0] dp2_ds0_out_mscbus;
wire     [31:0] dp2_ds1_out_mscbus;
wire     [31:0] dp2_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp2_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp2_gpio_out_2_buf_mscbus;
wire     [31:0] dp2_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp2_in_function_en_out_mscbus;
wire     [31:0] dp2_in_termination_en_out_mscbus;
wire     [31:0] dp2_inena_out_mscbus;
wire     [31:0] dp2_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp2_mode0_out_mscbus;
wire     [31:0] dp2_mode1_out_mscbus;
wire    [255:0] dp2_pes_en_out_mscbus;
wire     [31:0] dp2_pes_in_en_out_mscbus;
wire     [63:0] dp2_pes_safeval_out_mscbus;
wire    [159:0] dp2_pinmux_muxsel_out_mscbus;
wire     [31:0] dp2_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp2_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp2_pull_en_out_mscbus;
wire     [31:0] dp2_pull_type_out_mscbus;
wire     [31:0] dp2_schmitt_out_mscbus;
wire     [31:0] dp2_slew_out_mscbus;
wire     [31:0] dp3_GP_DATA_IN_out_mscbus;
wire     [31:0] dp3_amsel_out_mscbus;
wire     [31:0] dp3_async_in_from_pad_mscbus;
wire     [31:0] dp3_data_out_2_pinmux_mscbus;
wire     [31:0] dp3_dir_out_mscbus;
wire     [31:0] dp3_ds0_out_mscbus;
wire     [31:0] dp3_ds1_out_mscbus;
wire     [31:0] dp3_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp3_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp3_gpio_out_2_buf_mscbus;
wire     [31:0] dp3_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp3_in_function_en_out_mscbus;
wire     [31:0] dp3_in_termination_en_out_mscbus;
wire     [31:0] dp3_inena_out_mscbus;
wire     [31:0] dp3_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp3_mode0_out_mscbus;
wire     [31:0] dp3_mode1_out_mscbus;
wire    [255:0] dp3_pes_en_out_mscbus;
wire     [31:0] dp3_pes_in_en_out_mscbus;
wire     [63:0] dp3_pes_safeval_out_mscbus;
wire    [159:0] dp3_pinmux_muxsel_out_mscbus;
wire     [31:0] dp3_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp3_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp3_pull_en_out_mscbus;
wire     [31:0] dp3_pull_type_out_mscbus;
wire     [31:0] dp3_schmitt_out_mscbus;
wire     [31:0] dp3_slew_out_mscbus;
wire     [31:0] dp4_GP_DATA_IN_out_mscbus;
wire     [31:0] dp4_amsel_out_mscbus;
wire     [31:0] dp4_async_in_from_pad_mscbus;
wire     [31:0] dp4_data_out_2_pinmux_mscbus;
wire     [31:0] dp4_dir_out_mscbus;
wire     [31:0] dp4_ds0_out_mscbus;
wire     [31:0] dp4_ds1_out_mscbus;
wire     [31:0] dp4_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp4_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp4_gpio_out_2_buf_mscbus;
wire     [31:0] dp4_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp4_in_function_en_out_mscbus;
wire     [31:0] dp4_in_termination_en_out_mscbus;
wire     [31:0] dp4_inena_out_mscbus;
wire     [31:0] dp4_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp4_mode0_out_mscbus;
wire     [31:0] dp4_mode1_out_mscbus;
wire    [255:0] dp4_pes_en_out_mscbus;
wire     [31:0] dp4_pes_in_en_out_mscbus;
wire     [63:0] dp4_pes_safeval_out_mscbus;
wire    [159:0] dp4_pinmux_muxsel_out_mscbus;
wire     [31:0] dp4_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp4_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp4_pull_en_out_mscbus;
wire     [31:0] dp4_pull_type_out_mscbus;
wire     [31:0] dp4_schmitt_out_mscbus;
wire     [31:0] dp4_slew_out_mscbus;
wire     [31:0] dp5_GP_DATA_IN_out_mscbus;
wire     [31:0] dp5_amsel_out_mscbus;
wire     [31:0] dp5_async_in_from_pad_mscbus;
wire     [31:0] dp5_data_out_2_pinmux_mscbus;
wire     [31:0] dp5_dir_out_mscbus;
wire     [31:0] dp5_ds0_out_mscbus;
wire     [31:0] dp5_ds1_out_mscbus;
wire     [31:0] dp5_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp5_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp5_gpio_out_2_buf_mscbus;
wire     [31:0] dp5_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp5_in_function_en_out_mscbus;
wire     [31:0] dp5_in_termination_en_out_mscbus;
wire     [31:0] dp5_inena_out_mscbus;
wire     [31:0] dp5_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp5_mode0_out_mscbus;
wire     [31:0] dp5_mode1_out_mscbus;
wire    [255:0] dp5_pes_en_out_mscbus;
wire     [31:0] dp5_pes_in_en_out_mscbus;
wire     [63:0] dp5_pes_safeval_out_mscbus;
wire    [159:0] dp5_pinmux_muxsel_out_mscbus;
wire     [31:0] dp5_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp5_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp5_pull_en_out_mscbus;
wire     [31:0] dp5_pull_type_out_mscbus;
wire     [31:0] dp5_schmitt_out_mscbus;
wire     [31:0] dp5_slew_out_mscbus;
wire     [31:0] dp6_GP_DATA_IN_out_mscbus;
wire     [31:0] dp6_amsel_out_mscbus;
wire     [31:0] dp6_async_in_from_pad_mscbus;
wire     [31:0] dp6_data_out_2_pinmux_mscbus;
wire     [31:0] dp6_dir_out_mscbus;
wire     [31:0] dp6_ds0_out_mscbus;
wire     [31:0] dp6_ds1_out_mscbus;
wire     [31:0] dp6_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp6_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp6_gpio_out_2_buf_mscbus;
wire     [31:0] dp6_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp6_in_function_en_out_mscbus;
wire     [31:0] dp6_in_termination_en_out_mscbus;
wire     [31:0] dp6_inena_out_mscbus;
wire     [31:0] dp6_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp6_mode0_out_mscbus;
wire     [31:0] dp6_mode1_out_mscbus;
wire    [255:0] dp6_pes_en_out_mscbus;
wire     [31:0] dp6_pes_in_en_out_mscbus;
wire     [63:0] dp6_pes_safeval_out_mscbus;
wire    [159:0] dp6_pinmux_muxsel_out_mscbus;
wire     [31:0] dp6_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp6_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp6_pull_en_out_mscbus;
wire     [31:0] dp6_pull_type_out_mscbus;
wire     [31:0] dp6_schmitt_out_mscbus;
wire     [31:0] dp6_slew_out_mscbus;
wire     [31:0] dp7_GP_DATA_IN_out_mscbus;
wire     [31:0] dp7_amsel_out_mscbus;
wire     [31:0] dp7_async_in_from_pad_mscbus;
wire     [31:0] dp7_data_out_2_pinmux_mscbus;
wire     [31:0] dp7_dir_out_mscbus;
wire     [31:0] dp7_ds0_out_mscbus;
wire     [31:0] dp7_ds1_out_mscbus;
wire     [31:0] dp7_glitch_filter_bypass_out_mscbus;
wire     [63:0] dp7_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] dp7_gpio_out_2_buf_mscbus;
wire     [31:0] dp7_gpio_out_en_2_buf_mscbus;
wire   [1023:0] dp7_in_function_en_out_mscbus;
wire     [31:0] dp7_in_termination_en_out_mscbus;
wire     [31:0] dp7_inena_out_mscbus;
wire     [31:0] dp7_lvds_en_ctrl_out_mscbus;
wire     [31:0] dp7_mode0_out_mscbus;
wire     [31:0] dp7_mode1_out_mscbus;
wire    [255:0] dp7_pes_en_out_mscbus;
wire     [31:0] dp7_pes_in_en_out_mscbus;
wire     [63:0] dp7_pes_safeval_out_mscbus;
wire    [159:0] dp7_pinmux_muxsel_out_mscbus;
wire     [31:0] dp7_pinmuxdata_2_gpio_mscbus;
wire     [31:0] dp7_pinmuxen_2_gpio_mscbus;
wire     [31:0] dp7_pull_en_out_mscbus;
wire     [31:0] dp7_pull_type_out_mscbus;
wire     [31:0] dp7_schmitt_out_mscbus;
wire     [31:0] dp7_slew_out_mscbus;
wire     [31:0] mp0_GP_DATA_IN_out_mscbus;
wire     [31:0] mp0_amsel_out_mscbus;
wire     [31:0] mp0_async_in_from_pad_mscbus;
wire     [31:0] mp0_data_out_2_pinmux_mscbus;
wire     [31:0] mp0_dir_out_mscbus;
wire     [31:0] mp0_ds0_out_mscbus;
wire     [31:0] mp0_ds1_out_mscbus;
wire     [31:0] mp0_glitch_filter_bypass_out_mscbus;
wire     [63:0] mp0_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] mp0_gpio_out_2_buf_mscbus;
wire     [31:0] mp0_gpio_out_en_2_buf_mscbus;
wire   [1023:0] mp0_in_function_en_out_mscbus;
wire     [31:0] mp0_in_termination_en_out_mscbus;
wire     [31:0] mp0_inena_out_mscbus;
wire     [31:0] mp0_lvds_en_ctrl_out_mscbus;
wire     [31:0] mp0_mode0_out_mscbus;
wire     [31:0] mp0_mode1_out_mscbus;
wire    [255:0] mp0_pes_en_out_mscbus;
wire     [31:0] mp0_pes_in_en_out_mscbus;
wire     [63:0] mp0_pes_safeval_out_mscbus;
wire    [159:0] mp0_pinmux_muxsel_out_mscbus;
wire     [31:0] mp0_pinmuxdata_2_gpio_mscbus;
wire     [31:0] mp0_pinmuxen_2_gpio_mscbus;
wire     [31:0] mp0_pull_en_out_mscbus;
wire     [31:0] mp0_pull_type_out_mscbus;
wire     [31:0] mp0_schmitt_out_mscbus;
wire     [31:0] mp0_slew_out_mscbus;
wire     [31:0] mp1_GP_DATA_IN_out_mscbus;
wire     [31:0] mp1_amsel_out_mscbus;
wire     [31:0] mp1_async_in_from_pad_mscbus;
wire     [31:0] mp1_data_out_2_pinmux_mscbus;
wire     [31:0] mp1_dir_out_mscbus;
wire     [31:0] mp1_ds0_out_mscbus;
wire     [31:0] mp1_ds1_out_mscbus;
wire     [31:0] mp1_glitch_filter_bypass_out_mscbus;
wire     [63:0] mp1_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] mp1_gpio_out_2_buf_mscbus;
wire     [31:0] mp1_gpio_out_en_2_buf_mscbus;
wire   [1023:0] mp1_in_function_en_out_mscbus;
wire     [31:0] mp1_in_termination_en_out_mscbus;
wire     [31:0] mp1_inena_out_mscbus;
wire     [31:0] mp1_lvds_en_ctrl_out_mscbus;
wire     [31:0] mp1_mode0_out_mscbus;
wire     [31:0] mp1_mode1_out_mscbus;
wire    [255:0] mp1_pes_en_out_mscbus;
wire     [31:0] mp1_pes_in_en_out_mscbus;
wire     [63:0] mp1_pes_safeval_out_mscbus;
wire    [159:0] mp1_pinmux_muxsel_out_mscbus;
wire     [31:0] mp1_pinmuxdata_2_gpio_mscbus;
wire     [31:0] mp1_pinmuxen_2_gpio_mscbus;
wire     [31:0] mp1_pull_en_out_mscbus;
wire     [31:0] mp1_pull_type_out_mscbus;
wire     [31:0] mp1_schmitt_out_mscbus;
wire     [31:0] mp1_slew_out_mscbus;
wire     [31:0] mp2_GP_DATA_IN_out_mscbus;
wire     [31:0] mp2_amsel_out_mscbus;
wire     [31:0] mp2_async_in_from_pad_mscbus;
wire     [31:0] mp2_data_out_2_pinmux_mscbus;
wire     [31:0] mp2_dir_out_mscbus;
wire     [31:0] mp2_ds0_out_mscbus;
wire     [31:0] mp2_ds1_out_mscbus;
wire     [31:0] mp2_glitch_filter_bypass_out_mscbus;
wire     [63:0] mp2_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] mp2_gpio_out_2_buf_mscbus;
wire     [31:0] mp2_gpio_out_en_2_buf_mscbus;
wire   [1023:0] mp2_in_function_en_out_mscbus;
wire     [31:0] mp2_in_termination_en_out_mscbus;
wire     [31:0] mp2_inena_out_mscbus;
wire     [31:0] mp2_lvds_en_ctrl_out_mscbus;
wire     [31:0] mp2_mode0_out_mscbus;
wire     [31:0] mp2_mode1_out_mscbus;
wire    [255:0] mp2_pes_en_out_mscbus;
wire     [31:0] mp2_pes_in_en_out_mscbus;
wire     [63:0] mp2_pes_safeval_out_mscbus;
wire    [159:0] mp2_pinmux_muxsel_out_mscbus;
wire     [31:0] mp2_pinmuxdata_2_gpio_mscbus;
wire     [31:0] mp2_pinmuxen_2_gpio_mscbus;
wire     [31:0] mp2_pull_en_out_mscbus;
wire     [31:0] mp2_pull_type_out_mscbus;
wire     [31:0] mp2_schmitt_out_mscbus;
wire     [31:0] mp2_slew_out_mscbus;

// For DP ports (dp0 to dp7)
// MP Section (mp0 to mp2)
// AP Section (single instance)
pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(0)) I_b_DP0_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp0_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp0_inena_out_mscbus[0]),
  .dir_out_mscbus(dp0_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP0_0_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP0_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(1)) I_b_DP0_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp0_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp0_inena_out_mscbus[1]),
  .dir_out_mscbus(dp0_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_1_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(2)) I_b_DP0_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp0_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp0_inena_out_mscbus[2]),
  .dir_out_mscbus(dp0_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_2_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP0_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(3)) I_b_DP0_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp0_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp0_inena_out_mscbus[3]),
  .dir_out_mscbus(dp0_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_3_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_3_out_demux_peripheral_mscbus),
  .io_pad(DP0_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(4)) I_b_DP0_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp0_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp0_inena_out_mscbus[4]),
  .dir_out_mscbus(dp0_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_4_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP0_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(5)) I_b_DP0_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp0_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp0_inena_out_mscbus[5]),
  .dir_out_mscbus(dp0_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_5_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_5_out_demux_peripheral_mscbus),
  .io_pad(DP0_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(6)) I_b_DP0_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp0_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp0_inena_out_mscbus[6]),
  .dir_out_mscbus(dp0_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_6_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP0_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(7)) I_b_DP0_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp0_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp0_inena_out_mscbus[7]),
  .dir_out_mscbus(dp0_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_7_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_7_out_demux_peripheral_mscbus),
  .io_pad(DP0_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(8)) I_b_DP0_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp0_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp0_inena_out_mscbus[8]),
  .dir_out_mscbus(dp0_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_8_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_8_out_demux_peripheral_mscbus),
  .io_pad(DP0_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(9)) I_b_DP0_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp0_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp0_inena_out_mscbus[9]),
  .dir_out_mscbus(dp0_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_9_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_9_out_demux_peripheral_mscbus),
  .io_pad(DP0_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(10)) I_b_DP0_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp0_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp0_inena_out_mscbus[10]),
  .dir_out_mscbus(dp0_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_10_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP0_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(11)) I_b_DP0_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp0_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp0_inena_out_mscbus[11]),
  .dir_out_mscbus(dp0_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_11_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP0_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(12)) I_b_DP0_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp0_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp0_inena_out_mscbus[12]),
  .dir_out_mscbus(dp0_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_12_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP0_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(13)) I_b_DP0_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp0_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp0_inena_out_mscbus[13]),
  .dir_out_mscbus(dp0_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_13_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_13_out_demux_peripheral_mscbus),
  .io_pad(DP0_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(14)) I_b_DP0_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp0_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp0_inena_out_mscbus[14]),
  .dir_out_mscbus(dp0_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_14_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP0_14_out_demux_peripheral_mscbus),
  .io_pad(DP0_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(15)) I_b_DP0_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp0_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp0_inena_out_mscbus[15]),
  .dir_out_mscbus(dp0_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_15_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP0_15_out_demux_peripheral_mscbus),
  .io_pad(DP0_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(16)) I_b_DP0_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp0_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp0_inena_out_mscbus[16]),
  .dir_out_mscbus(dp0_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_16_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_16_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(17)) I_b_DP0_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp0_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp0_inena_out_mscbus[17]),
  .dir_out_mscbus(dp0_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_17_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_17_out_demux_peripheral_mscbus),
  .io_pad(DP0_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(18)) I_b_DP0_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp0_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp0_inena_out_mscbus[18]),
  .dir_out_mscbus(dp0_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_18_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_18_out_demux_peripheral_mscbus),
  .io_pad(DP0_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(19)) I_b_DP0_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp0_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp0_inena_out_mscbus[19]),
  .dir_out_mscbus(dp0_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_19_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP0_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(20)) I_b_DP0_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp0_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp0_inena_out_mscbus[20]),
  .dir_out_mscbus(dp0_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP0_20_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP0_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(21)) I_b_DP0_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp0_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp0_inena_out_mscbus[21]),
  .dir_out_mscbus(dp0_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_21_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_21_out_demux_peripheral_mscbus),
  .io_pad(DP0_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(22)) I_b_DP0_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp0_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp0_inena_out_mscbus[22]),
  .dir_out_mscbus(dp0_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_22_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_22_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(23)) I_b_DP0_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp0_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp0_inena_out_mscbus[23]),
  .dir_out_mscbus(dp0_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_23_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_23_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(24)) I_b_DP0_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp0_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp0_inena_out_mscbus[24]),
  .dir_out_mscbus(dp0_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_24_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_24_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(25)) I_b_DP0_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp0_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp0_inena_out_mscbus[25]),
  .dir_out_mscbus(dp0_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_25_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_25_out_demux_peripheral_mscbus),
  .io_pad(DP0_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(26)) I_b_DP0_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp0_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp0_inena_out_mscbus[26]),
  .dir_out_mscbus(dp0_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_26_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_26_out_demux_peripheral_mscbus),
  .io_pad(DP0_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(27)) I_b_DP0_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp0_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp0_inena_out_mscbus[27]),
  .dir_out_mscbus(dp0_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP0_27_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP0_27_out_demux_peripheral_mscbus),
  .io_pad(DP0_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(28)) I_b_DP0_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp0_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp0_inena_out_mscbus[28]),
  .dir_out_mscbus(dp0_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_28_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_28_out_demux_peripheral_mscbus),
  .io_pad(DP0_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(29)) I_b_DP0_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp0_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp0_inena_out_mscbus[29]),
  .dir_out_mscbus(dp0_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP0_29_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP0_29_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(30)) I_b_DP0_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp0_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp0_inena_out_mscbus[30]),
  .dir_out_mscbus(dp0_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP0_30_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP0_30_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP0_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(31)) I_b_DP0_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp0_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp0_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp0_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp0_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp0_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp0_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp0_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp0_inena_out_mscbus[31]),
  .dir_out_mscbus(dp0_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp0_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp0_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp0_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp0_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp0_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp0_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp0_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp0_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp0_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp0_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp0_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp0_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP0_31_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP0_31_out_demux_peripheral_mscbus),
  .io_pad(DP0_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(32)) I_b_DP1_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp1_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp1_inena_out_mscbus[0]),
  .dir_out_mscbus(dp1_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_0_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_0_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(33)) I_b_DP1_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp1_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp1_inena_out_mscbus[1]),
  .dir_out_mscbus(dp1_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_1_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(34)) I_b_DP1_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp1_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp1_inena_out_mscbus[2]),
  .dir_out_mscbus(dp1_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_2_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_2_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(35)) I_b_DP1_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp1_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp1_inena_out_mscbus[3]),
  .dir_out_mscbus(dp1_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_3_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_3_out_demux_peripheral_mscbus),
  .io_pad(DP1_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(36)) I_b_DP1_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp1_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp1_inena_out_mscbus[4]),
  .dir_out_mscbus(dp1_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_4_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_4_out_demux_peripheral_mscbus),
  .io_pad(DP1_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(37)) I_b_DP1_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp1_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp1_inena_out_mscbus[5]),
  .dir_out_mscbus(dp1_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_5_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_5_out_demux_peripheral_mscbus),
  .io_pad(DP1_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(38)) I_b_DP1_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp1_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp1_inena_out_mscbus[6]),
  .dir_out_mscbus(dp1_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_6_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_6_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(39)) I_b_DP1_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp1_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp1_inena_out_mscbus[7]),
  .dir_out_mscbus(dp1_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_7_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_7_out_demux_peripheral_mscbus),
  .io_pad(DP1_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(40)) I_b_DP1_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp1_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp1_inena_out_mscbus[8]),
  .dir_out_mscbus(dp1_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_8_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_8_out_demux_peripheral_mscbus),
  .io_pad(DP1_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(41)) I_b_DP1_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp1_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp1_inena_out_mscbus[9]),
  .dir_out_mscbus(dp1_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_9_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_9_out_demux_peripheral_mscbus),
  .io_pad(DP1_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(42)) I_b_DP1_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp1_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp1_inena_out_mscbus[10]),
  .dir_out_mscbus(dp1_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP1_10_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP1_10_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(43)) I_b_DP1_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp1_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp1_inena_out_mscbus[11]),
  .dir_out_mscbus(dp1_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP1_11_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP1_11_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(44)) I_b_DP1_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp1_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp1_inena_out_mscbus[12]),
  .dir_out_mscbus(dp1_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP1_12_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP1_12_out_demux_peripheral_mscbus),
  .io_pad(DP1_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(45)) I_b_DP1_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp1_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp1_inena_out_mscbus[13]),
  .dir_out_mscbus(dp1_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_13_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_13_out_demux_peripheral_mscbus),
  .io_pad(DP1_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(46)) I_b_DP1_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp1_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp1_inena_out_mscbus[14]),
  .dir_out_mscbus(dp1_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP1_14_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP1_14_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP1_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(47)) I_b_DP1_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp1_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp1_inena_out_mscbus[15]),
  .dir_out_mscbus(dp1_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_15_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_15_out_demux_peripheral_mscbus),
  .io_pad(DP1_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(48)) I_b_DP1_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp1_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp1_inena_out_mscbus[16]),
  .dir_out_mscbus(dp1_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_16_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_16_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(49)) I_b_DP1_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp1_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp1_inena_out_mscbus[17]),
  .dir_out_mscbus(dp1_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_17_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_17_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(50)) I_b_DP1_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp1_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp1_inena_out_mscbus[18]),
  .dir_out_mscbus(dp1_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_18_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_18_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(51)) I_b_DP1_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp1_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp1_inena_out_mscbus[19]),
  .dir_out_mscbus(dp1_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_19_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_19_out_demux_peripheral_mscbus),
  .io_pad(DP1_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(52)) I_b_DP1_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp1_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp1_inena_out_mscbus[20]),
  .dir_out_mscbus(dp1_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_20_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_20_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(53)) I_b_DP1_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp1_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp1_inena_out_mscbus[21]),
  .dir_out_mscbus(dp1_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_21_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_21_out_demux_peripheral_mscbus),
  .io_pad(DP1_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(54)) I_b_DP1_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp1_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp1_inena_out_mscbus[22]),
  .dir_out_mscbus(dp1_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_22_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_22_out_demux_peripheral_mscbus),
  .io_pad(DP1_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(55)) I_b_DP1_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp1_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp1_inena_out_mscbus[23]),
  .dir_out_mscbus(dp1_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_23_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_23_out_demux_peripheral_mscbus),
  .io_pad(DP1_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(56)) I_b_DP1_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp1_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp1_inena_out_mscbus[24]),
  .dir_out_mscbus(dp1_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_24_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_24_out_demux_peripheral_mscbus),
  .io_pad(DP1_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(57)) I_b_DP1_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp1_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp1_inena_out_mscbus[25]),
  .dir_out_mscbus(dp1_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP1_25_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP1_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(58)) I_b_DP1_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp1_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp1_inena_out_mscbus[26]),
  .dir_out_mscbus(dp1_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP1_26_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP1_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(59)) I_b_DP1_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp1_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp1_inena_out_mscbus[27]),
  .dir_out_mscbus(dp1_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP1_27_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP1_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(60)) I_b_DP1_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp1_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp1_inena_out_mscbus[28]),
  .dir_out_mscbus(dp1_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_28_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_28_out_demux_peripheral_mscbus),
  .io_pad(DP1_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(61)) I_b_DP1_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp1_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp1_inena_out_mscbus[29]),
  .dir_out_mscbus(dp1_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_29_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_29_out_demux_peripheral_mscbus),
  .io_pad(DP1_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(62)) I_b_DP1_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp1_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp1_inena_out_mscbus[30]),
  .dir_out_mscbus(dp1_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP1_30_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP1_30_out_demux_peripheral_mscbus),
  .io_pad(DP1_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(63)) I_b_DP1_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp1_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp1_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp1_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp1_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp1_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp1_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp1_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp1_inena_out_mscbus[31]),
  .dir_out_mscbus(dp1_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp1_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp1_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp1_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp1_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp1_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp1_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp1_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp1_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp1_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp1_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp1_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp1_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP1_31_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP1_31_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP1_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(64)) I_b_DP2_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp2_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp2_inena_out_mscbus[0]),
  .dir_out_mscbus(dp2_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_0_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_0_out_demux_peripheral_mscbus),
  .io_pad(DP2_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(65)) I_b_DP2_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp2_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp2_inena_out_mscbus[1]),
  .dir_out_mscbus(dp2_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_1_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(66)) I_b_DP2_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp2_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp2_inena_out_mscbus[2]),
  .dir_out_mscbus(dp2_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_2_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_2_out_demux_peripheral_mscbus),
  .io_pad(DP2_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(67)) I_b_DP2_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp2_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp2_inena_out_mscbus[3]),
  .dir_out_mscbus(dp2_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_3_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_3_out_demux_peripheral_mscbus),
  .io_pad(DP2_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(68)) I_b_DP2_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp2_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp2_inena_out_mscbus[4]),
  .dir_out_mscbus(dp2_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_4_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(69)) I_b_DP2_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp2_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp2_inena_out_mscbus[5]),
  .dir_out_mscbus(dp2_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_5_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(70)) I_b_DP2_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp2_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp2_inena_out_mscbus[6]),
  .dir_out_mscbus(dp2_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_6_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_6_out_demux_peripheral_mscbus),
  .io_pad(DP2_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(71)) I_b_DP2_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp2_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp2_inena_out_mscbus[7]),
  .dir_out_mscbus(dp2_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_7_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(72)) I_b_DP2_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp2_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp2_inena_out_mscbus[8]),
  .dir_out_mscbus(dp2_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_8_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(73)) I_b_DP2_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp2_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp2_inena_out_mscbus[9]),
  .dir_out_mscbus(dp2_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_9_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(74)) I_b_DP2_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp2_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp2_inena_out_mscbus[10]),
  .dir_out_mscbus(dp2_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_10_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(75)) I_b_DP2_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp2_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp2_inena_out_mscbus[11]),
  .dir_out_mscbus(dp2_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_11_in_mux_peripheral_mscbus[2:0]),
  .io_pad(DP2_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(76)) I_b_DP2_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp2_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp2_inena_out_mscbus[12]),
  .dir_out_mscbus(dp2_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_12_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_12_out_demux_peripheral_mscbus),
  .io_pad(DP2_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(77)) I_b_DP2_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp2_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp2_inena_out_mscbus[13]),
  .dir_out_mscbus(dp2_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_13_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_13_out_demux_peripheral_mscbus),
  .io_pad(DP2_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(78)) I_b_DP2_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp2_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp2_inena_out_mscbus[14]),
  .dir_out_mscbus(dp2_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_14_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(79)) I_b_DP2_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp2_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp2_inena_out_mscbus[15]),
  .dir_out_mscbus(dp2_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_15_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_15_out_demux_peripheral_mscbus),
  .io_pad(DP2_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(80)) I_b_DP2_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp2_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp2_inena_out_mscbus[16]),
  .dir_out_mscbus(dp2_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_16_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_16_out_demux_peripheral_mscbus),
  .io_pad(DP2_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(81)) I_b_DP2_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp2_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp2_inena_out_mscbus[17]),
  .dir_out_mscbus(dp2_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_17_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_17_out_demux_peripheral_mscbus),
  .io_pad(DP2_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(82)) I_b_DP2_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp2_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp2_inena_out_mscbus[18]),
  .dir_out_mscbus(dp2_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_18_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(83)) I_b_DP2_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp2_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp2_inena_out_mscbus[19]),
  .dir_out_mscbus(dp2_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_19_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP2_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(84)) I_b_DP2_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp2_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp2_inena_out_mscbus[20]),
  .dir_out_mscbus(dp2_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_20_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_20_out_demux_peripheral_mscbus),
  .io_pad(DP2_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(85)) I_b_DP2_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp2_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp2_inena_out_mscbus[21]),
  .dir_out_mscbus(dp2_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP2_21_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP2_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(86)) I_b_DP2_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp2_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp2_inena_out_mscbus[22]),
  .dir_out_mscbus(dp2_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP2_22_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP2_22_out_demux_peripheral_mscbus),
  .io_pad(DP2_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(87)) I_b_DP2_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp2_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp2_inena_out_mscbus[23]),
  .dir_out_mscbus(dp2_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP2_23_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP2_23_out_demux_peripheral_mscbus),
  .io_pad(DP2_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(88)) I_b_DP2_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp2_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp2_inena_out_mscbus[24]),
  .dir_out_mscbus(dp2_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP2_24_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP2_24_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP2_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(89)) I_b_DP2_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp2_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp2_inena_out_mscbus[25]),
  .dir_out_mscbus(dp2_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP2_25_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP2_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(90)) I_b_DP2_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp2_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp2_inena_out_mscbus[26]),
  .dir_out_mscbus(dp2_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_26_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_26_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP2_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(91)) I_b_DP2_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp2_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp2_inena_out_mscbus[27]),
  .dir_out_mscbus(dp2_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP2_27_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP2_27_out_demux_peripheral_mscbus),
  .io_pad(DP2_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(92)) I_b_DP2_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp2_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp2_inena_out_mscbus[28]),
  .dir_out_mscbus(dp2_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP2_28_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP2_28_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP2_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(93)) I_b_DP2_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp2_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp2_inena_out_mscbus[29]),
  .dir_out_mscbus(dp2_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP2_29_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP2_29_out_demux_peripheral_mscbus),
  .io_pad(DP2_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(94)) I_b_DP2_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp2_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp2_inena_out_mscbus[30]),
  .dir_out_mscbus(dp2_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP2_30_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP2_30_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP2_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(95)) I_b_DP2_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp2_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp2_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp2_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp2_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp2_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp2_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp2_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp2_inena_out_mscbus[31]),
  .dir_out_mscbus(dp2_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp2_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp2_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp2_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp0_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp2_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp2_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp2_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp2_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp2_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp2_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp2_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp2_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp2_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP2_31_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP2_31_out_demux_peripheral_mscbus),
  .io_pad(DP2_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(96)) I_b_DP3_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp3_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp3_inena_out_mscbus[0]),
  .dir_out_mscbus(dp3_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_0_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_0_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(97)) I_b_DP3_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp3_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp3_inena_out_mscbus[1]),
  .dir_out_mscbus(dp3_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_1_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(98)) I_b_DP3_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp3_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp3_inena_out_mscbus[2]),
  .dir_out_mscbus(dp3_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_2_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_2_out_demux_peripheral_mscbus),
  .io_pad(DP3_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(99)) I_b_DP3_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp3_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp3_inena_out_mscbus[3]),
  .dir_out_mscbus(dp3_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP3_3_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP3_3_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP3_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(100)) I_b_DP3_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp3_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp3_inena_out_mscbus[4]),
  .dir_out_mscbus(dp3_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_4_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_4_out_demux_peripheral_mscbus),
  .io_pad(DP3_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(101)) I_b_DP3_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp3_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp3_inena_out_mscbus[5]),
  .dir_out_mscbus(dp3_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_5_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_5_out_demux_peripheral_mscbus),
  .io_pad(DP3_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(102)) I_b_DP3_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp3_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp3_inena_out_mscbus[6]),
  .dir_out_mscbus(dp3_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_6_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_6_out_demux_peripheral_mscbus),
  .io_pad(DP3_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(103)) I_b_DP3_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp3_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp3_inena_out_mscbus[7]),
  .dir_out_mscbus(dp3_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_7_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_7_out_demux_peripheral_mscbus),
  .io_pad(DP3_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(104)) I_b_DP3_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp3_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp3_inena_out_mscbus[8]),
  .dir_out_mscbus(dp3_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_8_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_8_out_demux_peripheral_mscbus),
  .io_pad(DP3_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(105)) I_b_DP3_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp3_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp3_inena_out_mscbus[9]),
  .dir_out_mscbus(dp3_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_9_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_9_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(106)) I_b_DP3_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp3_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp3_inena_out_mscbus[10]),
  .dir_out_mscbus(dp3_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP3_10_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP3_10_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP3_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(107)) I_b_DP3_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp3_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp3_inena_out_mscbus[11]),
  .dir_out_mscbus(dp3_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_11_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_11_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(108)) I_b_DP3_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp3_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp3_inena_out_mscbus[12]),
  .dir_out_mscbus(dp3_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_12_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP3_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(109)) I_b_DP3_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp3_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp3_inena_out_mscbus[13]),
  .dir_out_mscbus(dp3_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_13_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_13_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(110)) I_b_DP3_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp3_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp3_inena_out_mscbus[14]),
  .dir_out_mscbus(dp3_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_14_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP3_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(111)) I_b_DP3_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp3_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp3_inena_out_mscbus[15]),
  .dir_out_mscbus(dp3_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_15_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_15_out_demux_peripheral_mscbus),
  .io_pad(DP3_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(112)) I_b_DP3_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp3_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp3_inena_out_mscbus[16]),
  .dir_out_mscbus(dp3_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_16_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_16_out_demux_peripheral_mscbus),
  .io_pad(DP3_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(113)) I_b_DP3_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp3_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp3_inena_out_mscbus[17]),
  .dir_out_mscbus(dp3_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP3_17_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP3_17_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(114)) I_b_DP3_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp3_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp3_inena_out_mscbus[18]),
  .dir_out_mscbus(dp3_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_18_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP3_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(115)) I_b_DP3_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp3_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp3_inena_out_mscbus[19]),
  .dir_out_mscbus(dp3_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_19_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP3_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(116)) I_b_DP3_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp3_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp3_inena_out_mscbus[20]),
  .dir_out_mscbus(dp3_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_20_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP3_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(117)) I_b_DP3_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp3_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp3_inena_out_mscbus[21]),
  .dir_out_mscbus(dp3_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP3_21_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP3_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(118)) I_b_DP3_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp3_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp3_inena_out_mscbus[22]),
  .dir_out_mscbus(dp3_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP3_22_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP3_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(119)) I_b_DP3_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp3_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp3_inena_out_mscbus[23]),
  .dir_out_mscbus(dp3_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP3_23_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP3_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(120)) I_b_DP3_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp3_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp3_inena_out_mscbus[24]),
  .dir_out_mscbus(dp3_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_24_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_24_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(121)) I_b_DP3_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp3_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp3_inena_out_mscbus[25]),
  .dir_out_mscbus(dp3_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP3_25_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP3_25_out_demux_peripheral_mscbus),
  .io_pad(DP3_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(122)) I_b_DP3_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp3_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp3_inena_out_mscbus[26]),
  .dir_out_mscbus(dp3_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_26_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_26_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(123)) I_b_DP3_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp3_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp3_inena_out_mscbus[27]),
  .dir_out_mscbus(dp3_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_27_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_27_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(124)) I_b_DP3_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp3_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp3_inena_out_mscbus[28]),
  .dir_out_mscbus(dp3_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_28_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_28_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP3_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(125)) I_b_DP3_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp3_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp3_inena_out_mscbus[29]),
  .dir_out_mscbus(dp3_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_29_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP3_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(126)) I_b_DP3_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp3_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp3_inena_out_mscbus[30]),
  .dir_out_mscbus(dp3_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP3_30_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP3_30_out_demux_peripheral_mscbus),
  .io_pad(DP3_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(127)) I_b_DP3_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp3_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp3_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp3_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp3_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp3_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp3_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp3_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp3_inena_out_mscbus[31]),
  .dir_out_mscbus(dp3_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp3_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp3_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp3_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp3_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp3_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp3_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp3_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp3_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp3_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp3_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp3_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp3_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp3_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP3_31_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP3_31_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP3_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(128)) I_b_DP4_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp4_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp4_inena_out_mscbus[0]),
  .dir_out_mscbus(dp4_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_0_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_0_out_demux_peripheral_mscbus),
  .io_pad(DP4_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(129)) I_b_DP4_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp4_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp4_inena_out_mscbus[1]),
  .dir_out_mscbus(dp4_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_1_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP4_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(130)) I_b_DP4_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp4_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp4_inena_out_mscbus[2]),
  .dir_out_mscbus(dp4_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_2_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_2_out_demux_peripheral_mscbus),
  .io_pad(DP4_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(131)) I_b_DP4_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp4_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp4_inena_out_mscbus[3]),
  .dir_out_mscbus(dp4_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_3_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_3_out_demux_peripheral_mscbus),
  .io_pad(DP4_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(132)) I_b_DP4_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp4_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp4_inena_out_mscbus[4]),
  .dir_out_mscbus(dp4_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_4_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP4_4_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(133)) I_b_DP4_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp4_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp4_inena_out_mscbus[5]),
  .dir_out_mscbus(dp4_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_5_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP4_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(134)) I_b_DP4_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp4_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp4_inena_out_mscbus[6]),
  .dir_out_mscbus(dp4_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP4_6_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP4_6_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(135)) I_b_DP4_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp4_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp4_inena_out_mscbus[7]),
  .dir_out_mscbus(dp4_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP4_7_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP4_7_out_demux_peripheral_mscbus),
  .io_pad(DP4_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(136)) I_b_DP4_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp4_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp4_inena_out_mscbus[8]),
  .dir_out_mscbus(dp4_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP4_8_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP4_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(137)) I_b_DP4_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp4_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp4_inena_out_mscbus[9]),
  .dir_out_mscbus(dp4_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_9_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_9_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(138)) I_b_DP4_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp4_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp4_inena_out_mscbus[10]),
  .dir_out_mscbus(dp4_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_10_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_10_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(139)) I_b_DP4_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp4_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp4_inena_out_mscbus[11]),
  .dir_out_mscbus(dp4_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP4_11_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP4_11_out_demux_peripheral_mscbus),
  .io_pad(DP4_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(140)) I_b_DP4_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp4_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp4_inena_out_mscbus[12]),
  .dir_out_mscbus(dp4_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_12_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_12_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(141)) I_b_DP4_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp4_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp4_inena_out_mscbus[13]),
  .dir_out_mscbus(dp4_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_13_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_13_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(142)) I_b_DP4_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp4_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp4_inena_out_mscbus[14]),
  .dir_out_mscbus(dp4_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_14_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_14_out_demux_peripheral_mscbus),
  .io_pad(DP4_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(143)) I_b_DP4_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp4_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp4_inena_out_mscbus[15]),
  .dir_out_mscbus(dp4_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_15_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_15_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP4_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(144)) I_b_DP4_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp4_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp4_inena_out_mscbus[16]),
  .dir_out_mscbus(dp4_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_16_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_16_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP4_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(145)) I_b_DP4_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp4_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp4_inena_out_mscbus[17]),
  .dir_out_mscbus(dp4_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_17_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_17_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP4_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(146)) I_b_DP4_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp4_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp4_inena_out_mscbus[18]),
  .dir_out_mscbus(dp4_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP4_18_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP4_18_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(147)) I_b_DP4_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp4_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp4_inena_out_mscbus[19]),
  .dir_out_mscbus(dp4_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_19_in_mux_peripheral_mscbus[2:0]),
  .io_pad(DP4_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(148)) I_b_DP4_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp4_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp4_inena_out_mscbus[20]),
  .dir_out_mscbus(dp4_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP4_20_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP4_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(149)) I_b_DP4_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp4_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp4_inena_out_mscbus[21]),
  .dir_out_mscbus(dp4_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP4_21_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP4_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(150)) I_b_DP4_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp4_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp4_inena_out_mscbus[22]),
  .dir_out_mscbus(dp4_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_22_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_22_out_demux_peripheral_mscbus),
  .io_pad(DP4_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(151)) I_b_DP4_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp4_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp4_inena_out_mscbus[23]),
  .dir_out_mscbus(dp4_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_23_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP4_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(152)) I_b_DP4_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp4_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp4_inena_out_mscbus[24]),
  .dir_out_mscbus(dp4_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_24_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP4_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(153)) I_b_DP4_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp4_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp4_inena_out_mscbus[25]),
  .dir_out_mscbus(dp4_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_25_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP4_25_out_demux_peripheral_mscbus),
  .io_pad(DP4_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(154)) I_b_DP4_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp4_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp4_inena_out_mscbus[26]),
  .dir_out_mscbus(dp4_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_26_in_mux_peripheral_mscbus[3:0]),
  .io_pad(DP4_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(155)) I_b_DP4_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp4_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp4_inena_out_mscbus[27]),
  .dir_out_mscbus(dp4_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_27_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_27_out_demux_peripheral_mscbus),
  .io_pad(DP4_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(156)) I_b_DP4_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp4_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp4_inena_out_mscbus[28]),
  .dir_out_mscbus(dp4_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP4_28_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP4_28_out_demux_peripheral_mscbus),
  .io_pad(DP4_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(157)) I_b_DP4_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp4_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp4_inena_out_mscbus[29]),
  .dir_out_mscbus(dp4_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_29_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP4_29_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(158)) I_b_DP4_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp4_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp4_inena_out_mscbus[30]),
  .dir_out_mscbus(dp4_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP4_30_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP4_30_out_demux_peripheral_mscbus),
  .io_pad(DP4_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(159)) I_b_DP4_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp4_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp4_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp4_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp4_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp4_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp4_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp4_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp4_inena_out_mscbus[31]),
  .dir_out_mscbus(dp4_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp4_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp4_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp4_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp4_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp4_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp4_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp4_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp4_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp4_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp4_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp4_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp4_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp4_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP4_31_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP4_31_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP4_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(160)) I_b_DP5_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp5_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp5_inena_out_mscbus[0]),
  .dir_out_mscbus(dp5_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP5_0_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP5_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(161)) I_b_DP5_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp5_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp5_inena_out_mscbus[1]),
  .dir_out_mscbus(dp5_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_1_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_1_out_demux_peripheral_mscbus),
  .io_pad(DP5_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(162)) I_b_DP5_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp5_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp5_inena_out_mscbus[2]),
  .dir_out_mscbus(dp5_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_2_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_2_out_demux_peripheral_mscbus),
  .io_pad(DP5_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(163)) I_b_DP5_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp5_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp5_inena_out_mscbus[3]),
  .dir_out_mscbus(dp5_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_3_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_3_out_demux_peripheral_mscbus),
  .io_pad(DP5_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(164)) I_b_DP5_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp5_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp5_inena_out_mscbus[4]),
  .dir_out_mscbus(dp5_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_4_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_4_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(165)) I_b_DP5_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp5_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp5_inena_out_mscbus[5]),
  .dir_out_mscbus(dp5_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_5_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_5_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(166)) I_b_DP5_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp5_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp5_inena_out_mscbus[6]),
  .dir_out_mscbus(dp5_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP5_6_in_mux_peripheral_mscbus[6:0]),
  .o_peripheral_in(DP5_6_out_demux_peripheral_mscbus),
  .io_pad(DP5_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(167)) I_b_DP5_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp5_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp5_inena_out_mscbus[7]),
  .dir_out_mscbus(dp5_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP5_7_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP5_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(168)) I_b_DP5_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp5_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp5_inena_out_mscbus[8]),
  .dir_out_mscbus(dp5_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP5_8_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP5_8_out_demux_peripheral_mscbus),
  .io_pad(DP5_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(4), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(169)) I_b_DP5_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp5_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp5_inena_out_mscbus[9]),
  .dir_out_mscbus(dp5_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP5_9_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP5_9_out_demux_peripheral_mscbus[3:0]),
  .io_pad(DP5_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(170)) I_b_DP5_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp5_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp5_inena_out_mscbus[10]),
  .dir_out_mscbus(dp5_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_10_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_10_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(171)) I_b_DP5_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp5_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp5_inena_out_mscbus[11]),
  .dir_out_mscbus(dp5_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP5_11_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP5_11_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP5_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(172)) I_b_DP5_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp5_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp5_inena_out_mscbus[12]),
  .dir_out_mscbus(dp5_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_12_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_12_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(173)) I_b_DP5_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp5_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp5_inena_out_mscbus[13]),
  .dir_out_mscbus(dp5_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_13_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_13_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(174)) I_b_DP5_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp5_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp5_inena_out_mscbus[14]),
  .dir_out_mscbus(dp5_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP5_14_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP5_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(175)) I_b_DP5_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp5_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp5_inena_out_mscbus[15]),
  .dir_out_mscbus(dp5_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_15_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_15_out_demux_peripheral_mscbus),
  .io_pad(DP5_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(176)) I_b_DP5_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp5_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp5_inena_out_mscbus[16]),
  .dir_out_mscbus(dp5_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_16_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_16_out_demux_peripheral_mscbus),
  .io_pad(DP5_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(177)) I_b_DP5_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp5_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp5_inena_out_mscbus[17]),
  .dir_out_mscbus(dp5_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_17_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_17_out_demux_peripheral_mscbus),
  .io_pad(DP5_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(178)) I_b_DP5_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp5_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp5_inena_out_mscbus[18]),
  .dir_out_mscbus(dp5_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_18_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP5_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(179)) I_b_DP5_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp5_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp5_inena_out_mscbus[19]),
  .dir_out_mscbus(dp5_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP5_19_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP5_19_out_demux_peripheral_mscbus),
  .io_pad(DP5_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(180)) I_b_DP5_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp5_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp5_inena_out_mscbus[20]),
  .dir_out_mscbus(dp5_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP5_20_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP5_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(181)) I_b_DP5_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp5_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp5_inena_out_mscbus[21]),
  .dir_out_mscbus(dp5_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_21_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_21_out_demux_peripheral_mscbus),
  .io_pad(DP5_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(182)) I_b_DP5_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp5_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp5_inena_out_mscbus[22]),
  .dir_out_mscbus(dp5_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP5_22_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP5_22_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(183)) I_b_DP5_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp5_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp5_inena_out_mscbus[23]),
  .dir_out_mscbus(dp5_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_23_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_23_out_demux_peripheral_mscbus),
  .io_pad(DP5_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(184)) I_b_DP5_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp5_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp5_inena_out_mscbus[24]),
  .dir_out_mscbus(dp5_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_24_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_24_out_demux_peripheral_mscbus),
  .io_pad(DP5_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(185)) I_b_DP5_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp5_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp5_inena_out_mscbus[25]),
  .dir_out_mscbus(dp5_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP5_25_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP5_25_out_demux_peripheral_mscbus),
  .io_pad(DP5_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(186)) I_b_DP5_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp5_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp5_inena_out_mscbus[26]),
  .dir_out_mscbus(dp5_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP5_26_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP5_26_out_demux_peripheral_mscbus),
  .io_pad(DP5_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(8), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(187)) I_b_DP5_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp5_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp5_inena_out_mscbus[27]),
  .dir_out_mscbus(dp5_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({8{1'b1}}),
  .i_peripheral_out(DP5_27_in_mux_peripheral_mscbus[7:0]),
  .io_pad(DP5_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(188)) I_b_DP5_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[28]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[28]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[28]),
  .slew_out_mscbus(dp5_slew_out_mscbus[28]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[28]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[28]),
  .inena_out_mscbus(dp5_inena_out_mscbus[28]),
  .dir_out_mscbus(dp5_dir_out_mscbus[28]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP5_28_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP5_28_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP5_28_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(189)) I_b_DP5_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[29]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[29]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[29]),
  .slew_out_mscbus(dp5_slew_out_mscbus[29]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[29]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[29]),
  .inena_out_mscbus(dp5_inena_out_mscbus[29]),
  .dir_out_mscbus(dp5_dir_out_mscbus[29]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[29]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP5_29_in_mux_peripheral_mscbus[6:0]),
  .o_peripheral_in(DP5_29_out_demux_peripheral_mscbus),
  .io_pad(DP5_29_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(190)) I_b_DP5_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[30]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[30]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[30]),
  .slew_out_mscbus(dp5_slew_out_mscbus[30]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[30]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[30]),
  .inena_out_mscbus(dp5_inena_out_mscbus[30]),
  .dir_out_mscbus(dp5_dir_out_mscbus[30]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP5_30_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP5_30_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP5_30_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(191)) I_b_DP5_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp5_amsel_out_mscbus[31]),
  .ds0_out_mscbus(dp5_ds0_out_mscbus[31]),
  .ds1_out_mscbus(dp5_ds1_out_mscbus[31]),
  .slew_out_mscbus(dp5_slew_out_mscbus[31]),
  .schmitt_out_mscbus(dp5_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(dp5_mode0_out_mscbus[31]),
  .mode1_out_mscbus(dp5_mode1_out_mscbus[31]),
  .inena_out_mscbus(dp5_inena_out_mscbus[31]),
  .dir_out_mscbus(dp5_dir_out_mscbus[31]),
  .pull_en_out_mscbus(dp5_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(dp5_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(dp5_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(dp5_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(dp5_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(dp5_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(dp5_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(dp5_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(dp5_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(dp5_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(dp5_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(dp5_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(dp5_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP5_31_in_mux_peripheral_mscbus[6:0]),
  .o_peripheral_in(DP5_31_out_demux_peripheral_mscbus),
  .io_pad(DP5_31_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(192)) I_b_DP6_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp6_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp6_inena_out_mscbus[0]),
  .dir_out_mscbus(dp6_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_0_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_0_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP6_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(193)) I_b_DP6_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp6_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp6_inena_out_mscbus[1]),
  .dir_out_mscbus(dp6_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_1_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(194)) I_b_DP6_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp6_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp6_inena_out_mscbus[2]),
  .dir_out_mscbus(dp6_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_2_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_2_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP6_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(195)) I_b_DP6_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp6_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp6_inena_out_mscbus[3]),
  .dir_out_mscbus(dp6_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP6_3_in_mux_peripheral_mscbus[6:0]),
  .o_peripheral_in(DP6_3_out_demux_peripheral_mscbus),
  .io_pad(DP6_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(196)) I_b_DP6_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp6_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp6_inena_out_mscbus[4]),
  .dir_out_mscbus(dp6_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_4_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_4_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(197)) I_b_DP6_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp6_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp6_inena_out_mscbus[5]),
  .dir_out_mscbus(dp6_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_5_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_5_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(198)) I_b_DP6_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp6_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp6_inena_out_mscbus[6]),
  .dir_out_mscbus(dp6_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_6_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_6_out_demux_peripheral_mscbus),
  .io_pad(DP6_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(199)) I_b_DP6_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp6_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp6_inena_out_mscbus[7]),
  .dir_out_mscbus(dp6_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_7_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_7_out_demux_peripheral_mscbus),
  .io_pad(DP6_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(200)) I_b_DP6_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp6_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp6_inena_out_mscbus[8]),
  .dir_out_mscbus(dp6_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP6_8_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP6_8_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(201)) I_b_DP6_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp6_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp6_inena_out_mscbus[9]),
  .dir_out_mscbus(dp6_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_9_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_9_out_demux_peripheral_mscbus),
  .io_pad(DP6_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(202)) I_b_DP6_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp6_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp6_inena_out_mscbus[10]),
  .dir_out_mscbus(dp6_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_10_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_10_out_demux_peripheral_mscbus),
  .io_pad(DP6_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(203)) I_b_DP6_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp6_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp6_inena_out_mscbus[11]),
  .dir_out_mscbus(dp6_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_11_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP6_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(204)) I_b_DP6_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp6_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp6_inena_out_mscbus[12]),
  .dir_out_mscbus(dp6_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_12_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_12_out_demux_peripheral_mscbus),
  .io_pad(DP6_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(205)) I_b_DP6_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp6_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp6_inena_out_mscbus[13]),
  .dir_out_mscbus(dp6_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_13_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_13_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(206)) I_b_DP6_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp6_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp6_inena_out_mscbus[14]),
  .dir_out_mscbus(dp6_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_14_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_14_out_demux_peripheral_mscbus),
  .io_pad(DP6_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(207)) I_b_DP6_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp6_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp6_inena_out_mscbus[15]),
  .dir_out_mscbus(dp6_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_15_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_15_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_15_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(208)) I_b_DP6_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[16]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[16]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[16]),
  .slew_out_mscbus(dp6_slew_out_mscbus[16]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[16]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[16]),
  .inena_out_mscbus(dp6_inena_out_mscbus[16]),
  .dir_out_mscbus(dp6_dir_out_mscbus[16]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_16_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_16_out_demux_peripheral_mscbus),
  .io_pad(DP6_16_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(209)) I_b_DP6_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[17]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[17]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[17]),
  .slew_out_mscbus(dp6_slew_out_mscbus[17]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[17]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[17]),
  .inena_out_mscbus(dp6_inena_out_mscbus[17]),
  .dir_out_mscbus(dp6_dir_out_mscbus[17]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[17]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP6_17_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP6_17_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(210)) I_b_DP6_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[18]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[18]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[18]),
  .slew_out_mscbus(dp6_slew_out_mscbus[18]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[18]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[18]),
  .inena_out_mscbus(dp6_inena_out_mscbus[18]),
  .dir_out_mscbus(dp6_dir_out_mscbus[18]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP6_18_in_mux_peripheral_mscbus[6:0]),
  .o_peripheral_in(DP6_18_out_demux_peripheral_mscbus),
  .io_pad(DP6_18_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(211)) I_b_DP6_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[19]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[19]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[19]),
  .slew_out_mscbus(dp6_slew_out_mscbus[19]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[19]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[19]),
  .inena_out_mscbus(dp6_inena_out_mscbus[19]),
  .dir_out_mscbus(dp6_dir_out_mscbus[19]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_19_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_19_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_19_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(7), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(212)) I_b_DP6_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[20]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[20]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[20]),
  .slew_out_mscbus(dp6_slew_out_mscbus[20]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[20]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[20]),
  .inena_out_mscbus(dp6_inena_out_mscbus[20]),
  .dir_out_mscbus(dp6_dir_out_mscbus[20]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({7{1'b1}}),
  .i_peripheral_out(DP6_20_in_mux_peripheral_mscbus[6:0]),
  .io_pad(DP6_20_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(213)) I_b_DP6_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[21]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[21]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[21]),
  .slew_out_mscbus(dp6_slew_out_mscbus[21]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[21]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[21]),
  .inena_out_mscbus(dp6_inena_out_mscbus[21]),
  .dir_out_mscbus(dp6_dir_out_mscbus[21]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP6_21_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP6_21_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP6_21_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(214)) I_b_DP6_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[22]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[22]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[22]),
  .slew_out_mscbus(dp6_slew_out_mscbus[22]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[22]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[22]),
  .inena_out_mscbus(dp6_inena_out_mscbus[22]),
  .dir_out_mscbus(dp6_dir_out_mscbus[22]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_22_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_22_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_22_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(215)) I_b_DP6_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[23]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[23]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[23]),
  .slew_out_mscbus(dp6_slew_out_mscbus[23]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[23]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[23]),
  .inena_out_mscbus(dp6_inena_out_mscbus[23]),
  .dir_out_mscbus(dp6_dir_out_mscbus[23]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_23_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_23_out_demux_peripheral_mscbus),
  .io_pad(DP6_23_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(216)) I_b_DP6_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[24]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[24]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[24]),
  .slew_out_mscbus(dp6_slew_out_mscbus[24]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[24]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[24]),
  .inena_out_mscbus(dp6_inena_out_mscbus[24]),
  .dir_out_mscbus(dp6_dir_out_mscbus[24]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP6_24_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP6_24_out_demux_peripheral_mscbus),
  .io_pad(DP6_24_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(217)) I_b_DP6_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[25]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[25]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[25]),
  .slew_out_mscbus(dp6_slew_out_mscbus[25]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[25]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[25]),
  .inena_out_mscbus(dp6_inena_out_mscbus[25]),
  .dir_out_mscbus(dp6_dir_out_mscbus[25]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[25]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_25_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP6_25_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP6_25_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(218)) I_b_DP6_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[26]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[26]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[26]),
  .slew_out_mscbus(dp6_slew_out_mscbus[26]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[26]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[26]),
  .inena_out_mscbus(dp6_inena_out_mscbus[26]),
  .dir_out_mscbus(dp6_dir_out_mscbus[26]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP6_26_in_mux_peripheral_mscbus[4:0]),
  .io_pad(DP6_26_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(219)) I_b_DP6_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp6_amsel_out_mscbus[27]),
  .ds0_out_mscbus(dp6_ds0_out_mscbus[27]),
  .ds1_out_mscbus(dp6_ds1_out_mscbus[27]),
  .slew_out_mscbus(dp6_slew_out_mscbus[27]),
  .schmitt_out_mscbus(dp6_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(dp6_mode0_out_mscbus[27]),
  .mode1_out_mscbus(dp6_mode1_out_mscbus[27]),
  .inena_out_mscbus(dp6_inena_out_mscbus[27]),
  .dir_out_mscbus(dp6_dir_out_mscbus[27]),
  .pull_en_out_mscbus(dp6_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(dp6_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(dp6_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(dp6_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(dp6_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(dp6_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(dp6_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(dp6_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(dp6_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(dp6_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(dp6_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(dp6_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(dp6_in_termination_en_out_mscbus[27]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP6_27_in_mux_peripheral_mscbus[2:0]),
  .io_pad(DP6_27_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(220)) I_b_DP7_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[0]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[0]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[0]),
  .slew_out_mscbus(dp7_slew_out_mscbus[0]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[0]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[0]),
  .inena_out_mscbus(dp7_inena_out_mscbus[0]),
  .dir_out_mscbus(dp7_dir_out_mscbus[0]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_0_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP7_0_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(221)) I_b_DP7_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[1]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[1]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[1]),
  .slew_out_mscbus(dp7_slew_out_mscbus[1]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[1]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[1]),
  .inena_out_mscbus(dp7_inena_out_mscbus[1]),
  .dir_out_mscbus(dp7_dir_out_mscbus[1]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(DP7_1_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(DP7_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP7_1_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(222)) I_b_DP7_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[2]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[2]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[2]),
  .slew_out_mscbus(dp7_slew_out_mscbus[2]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[2]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[2]),
  .inena_out_mscbus(dp7_inena_out_mscbus[2]),
  .dir_out_mscbus(dp7_dir_out_mscbus[2]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_2_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP7_2_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(223)) I_b_DP7_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[3]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[3]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[3]),
  .slew_out_mscbus(dp7_slew_out_mscbus[3]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[3]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[3]),
  .inena_out_mscbus(dp7_inena_out_mscbus[3]),
  .dir_out_mscbus(dp7_dir_out_mscbus[3]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_3_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP7_3_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(224)) I_b_DP7_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[4]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[4]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[4]),
  .slew_out_mscbus(dp7_slew_out_mscbus[4]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[4]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[4]),
  .inena_out_mscbus(dp7_inena_out_mscbus[4]),
  .dir_out_mscbus(dp7_dir_out_mscbus[4]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_4_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP7_4_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(225)) I_b_DP7_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[5]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[5]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[5]),
  .slew_out_mscbus(dp7_slew_out_mscbus[5]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[5]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[5]),
  .inena_out_mscbus(dp7_inena_out_mscbus[5]),
  .dir_out_mscbus(dp7_dir_out_mscbus[5]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_5_in_mux_peripheral_mscbus[5:0]),
  .io_pad(DP7_5_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(226)) I_b_DP7_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[6]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[6]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[6]),
  .slew_out_mscbus(dp7_slew_out_mscbus[6]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[6]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[6]),
  .inena_out_mscbus(dp7_inena_out_mscbus[6]),
  .dir_out_mscbus(dp7_dir_out_mscbus[6]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP7_6_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP7_6_out_demux_peripheral_mscbus),
  .io_pad(DP7_6_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(227)) I_b_DP7_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[7]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[7]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[7]),
  .slew_out_mscbus(dp7_slew_out_mscbus[7]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[7]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[7]),
  .inena_out_mscbus(dp7_inena_out_mscbus[7]),
  .dir_out_mscbus(dp7_dir_out_mscbus[7]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP7_7_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP7_7_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP7_7_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(6), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(228)) I_b_DP7_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[8]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[8]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[8]),
  .slew_out_mscbus(dp7_slew_out_mscbus[8]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[8]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[8]),
  .inena_out_mscbus(dp7_inena_out_mscbus[8]),
  .dir_out_mscbus(dp7_dir_out_mscbus[8]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({6{1'b1}}),
  .i_peripheral_out(DP7_8_in_mux_peripheral_mscbus[5:0]),
  .o_peripheral_in(DP7_8_out_demux_peripheral_mscbus),
  .io_pad(DP7_8_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(5), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(229)) I_b_DP7_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[9]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[9]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[9]),
  .slew_out_mscbus(dp7_slew_out_mscbus[9]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[9]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[9]),
  .inena_out_mscbus(dp7_inena_out_mscbus[9]),
  .dir_out_mscbus(dp7_dir_out_mscbus[9]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe({5{1'b1}}),
  .i_peripheral_out(DP7_9_in_mux_peripheral_mscbus[4:0]),
  .o_peripheral_in(DP7_9_out_demux_peripheral_mscbus),
  .io_pad(DP7_9_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(230)) I_b_DP7_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[10]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[10]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[10]),
  .slew_out_mscbus(dp7_slew_out_mscbus[10]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[10]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[10]),
  .inena_out_mscbus(dp7_inena_out_mscbus[10]),
  .dir_out_mscbus(dp7_dir_out_mscbus[10]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(DP7_10_in_mux_peripheral_mscbus),
  .o_peripheral_in(DP7_10_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP7_10_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(231)) I_b_DP7_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[11]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[11]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[11]),
  .slew_out_mscbus(dp7_slew_out_mscbus[11]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[11]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[11]),
  .inena_out_mscbus(dp7_inena_out_mscbus[11]),
  .dir_out_mscbus(dp7_dir_out_mscbus[11]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(DP7_11_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(DP7_11_out_demux_peripheral_mscbus),
  .io_pad(DP7_11_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(232)) I_b_DP7_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[12]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[12]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[12]),
  .slew_out_mscbus(dp7_slew_out_mscbus[12]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[12]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[12]),
  .inena_out_mscbus(dp7_inena_out_mscbus[12]),
  .dir_out_mscbus(dp7_dir_out_mscbus[12]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP7_12_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP7_12_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP7_12_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(233)) I_b_DP7_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[13]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[13]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[13]),
  .slew_out_mscbus(dp7_slew_out_mscbus[13]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[13]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[13]),
  .inena_out_mscbus(dp7_inena_out_mscbus[13]),
  .dir_out_mscbus(dp7_dir_out_mscbus[13]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(DP7_13_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(DP7_13_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP7_13_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(234)) I_b_DP7_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[14]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[14]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[14]),
  .slew_out_mscbus(dp7_slew_out_mscbus[14]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[14]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[14]),
  .inena_out_mscbus(dp7_inena_out_mscbus[14]),
  .dir_out_mscbus(dp7_dir_out_mscbus[14]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(DP7_14_in_mux_peripheral_mscbus),
  .o_peripheral_in(DP7_14_out_demux_peripheral_mscbus[2:0]),
  .io_pad(DP7_14_IO)
);

pinmux_with_io_dp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(235)) I_b_DP7_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(dp7_amsel_out_mscbus[15]),
  .ds0_out_mscbus(dp7_ds0_out_mscbus[15]),
  .ds1_out_mscbus(dp7_ds1_out_mscbus[15]),
  .slew_out_mscbus(dp7_slew_out_mscbus[15]),
  .schmitt_out_mscbus(dp7_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(dp7_mode0_out_mscbus[15]),
  .mode1_out_mscbus(dp7_mode1_out_mscbus[15]),
  .inena_out_mscbus(dp7_inena_out_mscbus[15]),
  .dir_out_mscbus(dp7_dir_out_mscbus[15]),
  .pull_en_out_mscbus(dp7_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(dp7_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(dp7_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(dp7_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(dp7_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(dp7_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(dp7_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(dp7_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(dp7_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(dp7_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(dp7_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(dp7_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(dp7_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(DP7_15_in_mux_peripheral_mscbus),
  .o_peripheral_in(DP7_15_out_demux_peripheral_mscbus[1:0]),
  .io_pad(DP7_15_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(236)) I_b_MP0_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[0]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[0]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[0]),
  .slew_out_mscbus(mp0_slew_out_mscbus[0]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[0]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[0]),
  .inena_out_mscbus(mp0_inena_out_mscbus[0]),
  .dir_out_mscbus(mp0_dir_out_mscbus[0]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_0_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_0_out_demux_peripheral_mscbus),
  .io_pad(MP0_0_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(237)) I_b_MP0_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[1]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[1]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[1]),
  .slew_out_mscbus(mp0_slew_out_mscbus[1]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[1]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[1]),
  .inena_out_mscbus(mp0_inena_out_mscbus[1]),
  .dir_out_mscbus(mp0_dir_out_mscbus[1]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_1_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_1_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_1_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(238)) I_b_MP0_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[2]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[2]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[2]),
  .slew_out_mscbus(mp0_slew_out_mscbus[2]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[2]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[2]),
  .inena_out_mscbus(mp0_inena_out_mscbus[2]),
  .dir_out_mscbus(mp0_dir_out_mscbus[2]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_2_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_2_out_demux_peripheral_mscbus),
  .io_pad(MP0_2_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(239)) I_b_MP0_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[3]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[3]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[3]),
  .slew_out_mscbus(mp0_slew_out_mscbus[3]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[3]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[3]),
  .inena_out_mscbus(mp0_inena_out_mscbus[3]),
  .dir_out_mscbus(mp0_dir_out_mscbus[3]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_3_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_3_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_3_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(240)) I_b_MP0_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[4]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[4]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[4]),
  .slew_out_mscbus(mp0_slew_out_mscbus[4]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[4]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[4]),
  .inena_out_mscbus(mp0_inena_out_mscbus[4]),
  .dir_out_mscbus(mp0_dir_out_mscbus[4]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_4_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_4_out_demux_peripheral_mscbus),
  .io_pad(MP0_4_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(241)) I_b_MP0_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[5]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[5]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[5]),
  .slew_out_mscbus(mp0_slew_out_mscbus[5]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[5]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[5]),
  .inena_out_mscbus(mp0_inena_out_mscbus[5]),
  .dir_out_mscbus(mp0_dir_out_mscbus[5]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[5]),
  .o_peripheral_in(MP0_5_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_5_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(242)) I_b_MP0_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[6]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[6]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[6]),
  .slew_out_mscbus(mp0_slew_out_mscbus[6]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[6]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[6]),
  .inena_out_mscbus(mp0_inena_out_mscbus[6]),
  .dir_out_mscbus(mp0_dir_out_mscbus[6]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_6_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_6_out_demux_peripheral_mscbus),
  .io_pad(MP0_6_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(243)) I_b_MP0_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[7]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[7]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[7]),
  .slew_out_mscbus(mp0_slew_out_mscbus[7]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[7]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[7]),
  .inena_out_mscbus(mp0_inena_out_mscbus[7]),
  .dir_out_mscbus(mp0_dir_out_mscbus[7]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_7_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_7_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_7_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(244)) I_b_MP0_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[8]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[8]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[8]),
  .slew_out_mscbus(mp0_slew_out_mscbus[8]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[8]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[8]),
  .inena_out_mscbus(mp0_inena_out_mscbus[8]),
  .dir_out_mscbus(mp0_dir_out_mscbus[8]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(MP0_8_in_mux_peripheral_mscbus[3:0]),
  .o_peripheral_in(MP0_8_out_demux_peripheral_mscbus),
  .io_pad(MP0_8_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(245)) I_b_MP0_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[9]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[9]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[9]),
  .slew_out_mscbus(mp0_slew_out_mscbus[9]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[9]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[9]),
  .inena_out_mscbus(mp0_inena_out_mscbus[9]),
  .dir_out_mscbus(mp0_dir_out_mscbus[9]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP0_9_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP0_9_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP0_9_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(246)) I_b_MP0_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[10]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[10]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[10]),
  .slew_out_mscbus(mp0_slew_out_mscbus[10]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[10]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[10]),
  .inena_out_mscbus(mp0_inena_out_mscbus[10]),
  .dir_out_mscbus(mp0_dir_out_mscbus[10]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_10_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_10_out_demux_peripheral_mscbus),
  .io_pad(MP0_10_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(247)) I_b_MP0_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[11]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[11]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[11]),
  .slew_out_mscbus(mp0_slew_out_mscbus[11]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[11]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[11]),
  .inena_out_mscbus(mp0_inena_out_mscbus[11]),
  .dir_out_mscbus(mp0_dir_out_mscbus[11]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[11]),
  .o_peripheral_in(MP0_11_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP0_11_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(248)) I_b_MP0_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[12]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[12]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[12]),
  .slew_out_mscbus(mp0_slew_out_mscbus[12]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[12]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[12]),
  .inena_out_mscbus(mp0_inena_out_mscbus[12]),
  .dir_out_mscbus(mp0_dir_out_mscbus[12]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_12_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP0_12_out_demux_peripheral_mscbus),
  .io_pad(MP0_12_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(249)) I_b_MP0_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[13]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[13]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[13]),
  .slew_out_mscbus(mp0_slew_out_mscbus[13]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[13]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[13]),
  .inena_out_mscbus(mp0_inena_out_mscbus[13]),
  .dir_out_mscbus(mp0_dir_out_mscbus[13]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP0_13_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP0_13_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP0_13_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(250)) I_b_MP0_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[14]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[14]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[14]),
  .slew_out_mscbus(mp0_slew_out_mscbus[14]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[14]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[14]),
  .inena_out_mscbus(mp0_inena_out_mscbus[14]),
  .dir_out_mscbus(mp0_dir_out_mscbus[14]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(MP0_14_in_mux_peripheral_mscbus[3:0]),
  .io_pad(MP0_14_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(251)) I_b_MP0_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[15]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[15]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[15]),
  .slew_out_mscbus(mp0_slew_out_mscbus[15]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[15]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[15]),
  .inena_out_mscbus(mp0_inena_out_mscbus[15]),
  .dir_out_mscbus(mp0_dir_out_mscbus[15]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_15_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_15_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_15_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(252)) I_b_MP0_16(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[16]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[16]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[16]),
  .slew_out_mscbus(mp0_slew_out_mscbus[16]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[16]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[16]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[16]),
  .inena_out_mscbus(mp0_inena_out_mscbus[16]),
  .dir_out_mscbus(mp0_dir_out_mscbus[16]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[16]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[16]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[84:80]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[543:512]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[16]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[16]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[16]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[16]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[16]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[16]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[16]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[16]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[16]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(MP0_16_in_mux_peripheral_mscbus[3:0]),
  .io_pad(MP0_16_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(253)) I_b_MP0_17(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[17]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[17]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[17]),
  .slew_out_mscbus(mp0_slew_out_mscbus[17]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[17]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[17]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[17]),
  .inena_out_mscbus(mp0_inena_out_mscbus[17]),
  .dir_out_mscbus(mp0_dir_out_mscbus[17]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[17]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[17]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[89:85]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[575:544]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[17]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[17]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[17]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[17]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[17]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[17]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[17]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[17]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[17]),
  .o_peripheral_in(MP0_17_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_17_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(254)) I_b_MP0_18(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[18]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[18]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[18]),
  .slew_out_mscbus(mp0_slew_out_mscbus[18]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[18]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[18]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[18]),
  .inena_out_mscbus(mp0_inena_out_mscbus[18]),
  .dir_out_mscbus(mp0_dir_out_mscbus[18]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[18]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[18]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[94:90]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[607:576]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[18]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[18]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[18]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[18]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[18]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[18]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[18]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[18]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[18]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(MP0_18_in_mux_peripheral_mscbus[3:0]),
  .io_pad(MP0_18_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(255)) I_b_MP0_19(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[19]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[19]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[19]),
  .slew_out_mscbus(mp0_slew_out_mscbus[19]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[19]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[19]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[19]),
  .inena_out_mscbus(mp0_inena_out_mscbus[19]),
  .dir_out_mscbus(mp0_dir_out_mscbus[19]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[19]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[19]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[99:95]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[639:608]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[19]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[19]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[19]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[19]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[19]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[19]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[19]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[19]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[19]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_19_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_19_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_19_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(4), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(256)) I_b_MP0_20(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[20]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[20]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[20]),
  .slew_out_mscbus(mp0_slew_out_mscbus[20]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[20]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[20]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[20]),
  .inena_out_mscbus(mp0_inena_out_mscbus[20]),
  .dir_out_mscbus(mp0_dir_out_mscbus[20]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[20]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[20]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[104:100]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[671:640]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[20]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[20]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[20]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[20]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[20]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[20]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[20]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[20]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[20]),
  .i_peripheral_oe({4{1'b1}}),
  .i_peripheral_out(MP0_20_in_mux_peripheral_mscbus[3:0]),
  .io_pad(MP0_20_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(257)) I_b_MP0_21(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[21]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[21]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[21]),
  .slew_out_mscbus(mp0_slew_out_mscbus[21]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[21]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[21]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[21]),
  .inena_out_mscbus(mp0_inena_out_mscbus[21]),
  .dir_out_mscbus(mp0_dir_out_mscbus[21]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[21]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[21]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[109:105]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[703:672]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[21]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[21]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[21]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[21]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[21]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[21]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[21]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[21]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[21]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_21_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_21_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_21_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(258)) I_b_MP0_22(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[22]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[22]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[22]),
  .slew_out_mscbus(mp0_slew_out_mscbus[22]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[22]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[22]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[22]),
  .inena_out_mscbus(mp0_inena_out_mscbus[22]),
  .dir_out_mscbus(mp0_dir_out_mscbus[22]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[22]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[22]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[114:110]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[735:704]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[22]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[22]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[22]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[22]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[22]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[22]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[22]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[22]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[22]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_22_in_mux_peripheral_mscbus[2:0]),
  .io_pad(MP0_22_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(259)) I_b_MP0_23(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[23]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[23]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[23]),
  .slew_out_mscbus(mp0_slew_out_mscbus[23]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[23]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[23]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[23]),
  .inena_out_mscbus(mp0_inena_out_mscbus[23]),
  .dir_out_mscbus(mp0_dir_out_mscbus[23]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[23]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[23]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[119:115]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[767:736]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[23]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[23]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[23]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[23]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[23]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[23]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[23]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[23]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[23]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP0_23_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP0_23_out_demux_peripheral_mscbus),
  .io_pad(MP0_23_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(260)) I_b_MP0_24(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[24]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[24]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[24]),
  .slew_out_mscbus(mp0_slew_out_mscbus[24]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[24]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[24]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[24]),
  .inena_out_mscbus(mp0_inena_out_mscbus[24]),
  .dir_out_mscbus(mp0_dir_out_mscbus[24]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[24]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[24]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[124:120]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[799:768]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[24]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[24]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[24]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[24]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[24]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[24]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[24]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[24]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[24]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP0_24_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP0_24_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_24_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(261)) I_b_MP0_25(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[25]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[25]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[25]),
  .slew_out_mscbus(mp0_slew_out_mscbus[25]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[25]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[25]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[25]),
  .inena_out_mscbus(mp0_inena_out_mscbus[25]),
  .dir_out_mscbus(mp0_dir_out_mscbus[25]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[25]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[25]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[129:125]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[831:800]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[25]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[25]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[25]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[25]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[25]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[25]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[25]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[25]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[25]),
  .o_peripheral_in(MP0_25_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP0_25_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(262)) I_b_MP0_26(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[26]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[26]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[26]),
  .slew_out_mscbus(mp0_slew_out_mscbus[26]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[26]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[26]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[26]),
  .inena_out_mscbus(mp0_inena_out_mscbus[26]),
  .dir_out_mscbus(mp0_dir_out_mscbus[26]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[26]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[26]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[134:130]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[863:832]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[26]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[26]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[26]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[26]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[26]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[26]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[26]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[26]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[26]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_26_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_26_out_demux_peripheral_mscbus),
  .io_pad(MP0_26_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(263)) I_b_MP0_27(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[27]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[27]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[27]),
  .slew_out_mscbus(mp0_slew_out_mscbus[27]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[27]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[27]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[27]),
  .inena_out_mscbus(mp0_inena_out_mscbus[27]),
  .dir_out_mscbus(mp0_dir_out_mscbus[27]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[27]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[27]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[139:135]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[895:864]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[27]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[27]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[27]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[27]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[27]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[27]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[27]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[27]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[27]),
  .o_peripheral_in(MP0_27_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP0_27_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(264)) I_b_MP0_28(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[28]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[28]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[28]),
  .slew_out_mscbus(mp0_slew_out_mscbus[28]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[28]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[28]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[28]),
  .inena_out_mscbus(mp0_inena_out_mscbus[28]),
  .dir_out_mscbus(mp0_dir_out_mscbus[28]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[28]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[28]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[144:140]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[927:896]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[28]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[28]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[28]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[28]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[28]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[28]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[28]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[28]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[28]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_28_in_mux_peripheral_mscbus[2:0]),
  .io_pad(MP0_28_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(265)) I_b_MP0_29(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[29]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[29]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[29]),
  .slew_out_mscbus(mp0_slew_out_mscbus[29]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[29]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[29]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[29]),
  .inena_out_mscbus(mp0_inena_out_mscbus[29]),
  .dir_out_mscbus(mp0_dir_out_mscbus[29]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[29]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[29]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[149:145]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[959:928]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[29]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[29]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[29]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[29]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[29]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[29]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[29]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[29]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[29]),
  .o_peripheral_in(MP0_29_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP0_29_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(266)) I_b_MP0_30(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[30]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[30]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[30]),
  .slew_out_mscbus(mp0_slew_out_mscbus[30]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[30]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[30]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[30]),
  .inena_out_mscbus(mp0_inena_out_mscbus[30]),
  .dir_out_mscbus(mp0_dir_out_mscbus[30]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[30]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[30]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[154:150]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[991:960]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[30]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[30]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[30]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[30]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[30]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[30]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[30]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[30]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[30]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP0_30_in_mux_peripheral_mscbus[2:0]),
  .io_pad(MP0_30_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(267)) I_b_MP0_31(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp0_amsel_out_mscbus[31]),
  .ds0_out_mscbus(mp0_ds0_out_mscbus[31]),
  .ds1_out_mscbus(mp0_ds1_out_mscbus[31]),
  .slew_out_mscbus(mp0_slew_out_mscbus[31]),
  .schmitt_out_mscbus(mp0_schmitt_out_mscbus[31]),
  .mode0_out_mscbus(mp0_mode0_out_mscbus[31]),
  .mode1_out_mscbus(mp0_mode1_out_mscbus[31]),
  .inena_out_mscbus(mp0_inena_out_mscbus[31]),
  .dir_out_mscbus(mp0_dir_out_mscbus[31]),
  .pull_en_out_mscbus(mp0_pull_en_out_mscbus[31]),
  .pull_type_out_mscbus(mp0_pull_type_out_mscbus[31]),
  .pinmux_muxsel_out_mscbus(mp0_pinmux_muxsel_out_mscbus[159:155]),
  .in_function_en_out_mscbus(mp0_in_function_en_out_mscbus[1023:992]),
  .async_in_from_pad_mscbus(mp0_async_in_from_pad_mscbus[31]),
  .gpio_out_2_buf_mscbus(mp0_gpio_out_2_buf_mscbus[31]),
  .gpio_out_en_2_buf_mscbus(mp0_gpio_out_en_2_buf_mscbus[31]),
  .pinmuxdata_2_gpio_mscbus(mp0_pinmuxdata_2_gpio_mscbus[31]),
  .pinmuxen_2_gpio_mscbus(mp0_pinmuxen_2_gpio_mscbus[31]),
  .GP_DATA_IN_out_mscbus(mp0_GP_DATA_IN_out_mscbus[31]),
  .data_out_2_pinmux_mscbus(mp0_data_out_2_pinmux_mscbus[31]),
  .lvds_en_ctrl_out_mscbus(mp0_lvds_en_ctrl_out_mscbus[31]),
  .in_termination_en_out_mscbus(mp0_in_termination_en_out_mscbus[31]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP0_31_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP0_31_out_demux_peripheral_mscbus),
  .io_pad(MP0_31_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(268)) I_b_MP1_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[0]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[0]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[0]),
  .slew_out_mscbus(mp1_slew_out_mscbus[0]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[0]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[0]),
  .inena_out_mscbus(mp1_inena_out_mscbus[0]),
  .dir_out_mscbus(mp1_dir_out_mscbus[0]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP1_0_in_mux_peripheral_mscbus[2:0]),
  .io_pad(MP1_0_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(269)) I_b_MP1_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[1]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[1]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[1]),
  .slew_out_mscbus(mp1_slew_out_mscbus[1]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[1]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[1]),
  .inena_out_mscbus(mp1_inena_out_mscbus[1]),
  .dir_out_mscbus(mp1_dir_out_mscbus[1]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP1_1_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP1_1_out_demux_peripheral_mscbus),
  .io_pad(MP1_1_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(270)) I_b_MP1_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[2]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[2]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[2]),
  .slew_out_mscbus(mp1_slew_out_mscbus[2]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[2]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[2]),
  .inena_out_mscbus(mp1_inena_out_mscbus[2]),
  .dir_out_mscbus(mp1_dir_out_mscbus[2]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP1_2_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP1_2_out_demux_peripheral_mscbus),
  .io_pad(MP1_2_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(0), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(271)) I_b_MP1_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[3]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[3]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[3]),
  .slew_out_mscbus(mp1_slew_out_mscbus[3]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[3]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[3]),
  .inena_out_mscbus(mp1_inena_out_mscbus[3]),
  .dir_out_mscbus(mp1_dir_out_mscbus[3]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[3]),
  .o_peripheral_in(MP1_3_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP1_3_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(272)) I_b_MP1_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[4]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[4]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[4]),
  .slew_out_mscbus(mp1_slew_out_mscbus[4]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[4]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[4]),
  .inena_out_mscbus(mp1_inena_out_mscbus[4]),
  .dir_out_mscbus(mp1_dir_out_mscbus[4]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_4_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_4_out_demux_peripheral_mscbus),
  .io_pad(MP1_4_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(273)) I_b_MP1_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[5]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[5]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[5]),
  .slew_out_mscbus(mp1_slew_out_mscbus[5]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[5]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[5]),
  .inena_out_mscbus(mp1_inena_out_mscbus[5]),
  .dir_out_mscbus(mp1_dir_out_mscbus[5]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_5_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_5_out_demux_peripheral_mscbus),
  .io_pad(MP1_5_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(274)) I_b_MP1_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[6]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[6]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[6]),
  .slew_out_mscbus(mp1_slew_out_mscbus[6]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[6]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[6]),
  .inena_out_mscbus(mp1_inena_out_mscbus[6]),
  .dir_out_mscbus(mp1_dir_out_mscbus[6]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_6_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_6_out_demux_peripheral_mscbus),
  .io_pad(MP1_6_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(275)) I_b_MP1_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[7]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[7]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[7]),
  .slew_out_mscbus(mp1_slew_out_mscbus[7]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[7]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[7]),
  .inena_out_mscbus(mp1_inena_out_mscbus[7]),
  .dir_out_mscbus(mp1_dir_out_mscbus[7]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_7_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_7_out_demux_peripheral_mscbus),
  .io_pad(MP1_7_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(276)) I_b_MP1_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[8]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[8]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[8]),
  .slew_out_mscbus(mp1_slew_out_mscbus[8]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[8]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[8]),
  .inena_out_mscbus(mp1_inena_out_mscbus[8]),
  .dir_out_mscbus(mp1_dir_out_mscbus[8]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_8_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_8_out_demux_peripheral_mscbus),
  .io_pad(MP1_8_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(277)) I_b_MP1_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[9]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[9]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[9]),
  .slew_out_mscbus(mp1_slew_out_mscbus[9]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[9]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[9]),
  .inena_out_mscbus(mp1_inena_out_mscbus[9]),
  .dir_out_mscbus(mp1_dir_out_mscbus[9]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_9_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP1_9_out_demux_peripheral_mscbus),
  .io_pad(MP1_9_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(278)) I_b_MP1_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[10]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[10]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[10]),
  .slew_out_mscbus(mp1_slew_out_mscbus[10]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[10]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[10]),
  .inena_out_mscbus(mp1_inena_out_mscbus[10]),
  .dir_out_mscbus(mp1_dir_out_mscbus[10]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP1_10_in_mux_peripheral_mscbus[1:0]),
  .io_pad(MP1_10_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(279)) I_b_MP1_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[11]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[11]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[11]),
  .slew_out_mscbus(mp1_slew_out_mscbus[11]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[11]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[11]),
  .inena_out_mscbus(mp1_inena_out_mscbus[11]),
  .dir_out_mscbus(mp1_dir_out_mscbus[11]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP1_11_in_mux_peripheral_mscbus[1:0]),
  .io_pad(MP1_11_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(280)) I_b_MP1_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[12]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[12]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[12]),
  .slew_out_mscbus(mp1_slew_out_mscbus[12]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[12]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[12]),
  .inena_out_mscbus(mp1_inena_out_mscbus[12]),
  .dir_out_mscbus(mp1_dir_out_mscbus[12]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_12_in_mux_peripheral_mscbus),
  .io_pad(MP1_12_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(281)) I_b_MP1_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[13]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[13]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[13]),
  .slew_out_mscbus(mp1_slew_out_mscbus[13]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[13]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[13]),
  .inena_out_mscbus(mp1_inena_out_mscbus[13]),
  .dir_out_mscbus(mp1_dir_out_mscbus[13]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_13_in_mux_peripheral_mscbus),
  .io_pad(MP1_13_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(282)) I_b_MP1_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[14]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[14]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[14]),
  .slew_out_mscbus(mp1_slew_out_mscbus[14]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[14]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[14]),
  .inena_out_mscbus(mp1_inena_out_mscbus[14]),
  .dir_out_mscbus(mp1_dir_out_mscbus[14]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_14_in_mux_peripheral_mscbus),
  .io_pad(MP1_14_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(0), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(283)) I_b_MP1_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp1_amsel_out_mscbus[15]),
  .ds0_out_mscbus(mp1_ds0_out_mscbus[15]),
  .ds1_out_mscbus(mp1_ds1_out_mscbus[15]),
  .slew_out_mscbus(mp1_slew_out_mscbus[15]),
  .schmitt_out_mscbus(mp1_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(mp1_mode0_out_mscbus[15]),
  .mode1_out_mscbus(mp1_mode1_out_mscbus[15]),
  .inena_out_mscbus(mp1_inena_out_mscbus[15]),
  .dir_out_mscbus(mp1_dir_out_mscbus[15]),
  .pull_en_out_mscbus(mp1_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(mp1_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(mp1_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(mp1_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(mp1_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(mp1_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(mp1_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(mp1_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(mp1_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(mp1_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(mp1_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(mp1_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(mp1_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP1_15_in_mux_peripheral_mscbus),
  .io_pad(MP1_15_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(284)) I_b_MP2_0(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[0]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[0]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[0]),
  .slew_out_mscbus(mp2_slew_out_mscbus[0]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[0]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[0]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[0]),
  .inena_out_mscbus(mp2_inena_out_mscbus[0]),
  .dir_out_mscbus(mp2_dir_out_mscbus[0]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[0]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[0]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[4:0]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[31:0]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[0]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[0]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[0]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[0]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[0]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[0]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[0]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[0]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[0]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_0_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_0_out_demux_peripheral_mscbus),
  .io_pad(MP2_0_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(285)) I_b_MP2_1(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[1]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[1]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[1]),
  .slew_out_mscbus(mp2_slew_out_mscbus[1]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[1]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[1]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[1]),
  .inena_out_mscbus(mp2_inena_out_mscbus[1]),
  .dir_out_mscbus(mp2_dir_out_mscbus[1]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[1]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[1]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[9:5]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[63:32]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[1]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[1]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[1]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[1]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[1]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[1]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[1]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[1]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[1]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP2_1_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP2_1_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP2_1_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(286)) I_b_MP2_2(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[2]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[2]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[2]),
  .slew_out_mscbus(mp2_slew_out_mscbus[2]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[2]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[2]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[2]),
  .inena_out_mscbus(mp2_inena_out_mscbus[2]),
  .dir_out_mscbus(mp2_dir_out_mscbus[2]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[2]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[2]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[14:10]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[95:64]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[2]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[2]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[2]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[2]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[2]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[2]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[2]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[2]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[2]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_2_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_2_out_demux_peripheral_mscbus),
  .io_pad(MP2_2_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(287)) I_b_MP2_3(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[3]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[3]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[3]),
  .slew_out_mscbus(mp2_slew_out_mscbus[3]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[3]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[3]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[3]),
  .inena_out_mscbus(mp2_inena_out_mscbus[3]),
  .dir_out_mscbus(mp2_dir_out_mscbus[3]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[3]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[3]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[19:15]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[127:96]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[3]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[3]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[3]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[3]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[3]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[3]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[3]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[3]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[3]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_3_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_3_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP2_3_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(288)) I_b_MP2_4(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[4]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[4]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[4]),
  .slew_out_mscbus(mp2_slew_out_mscbus[4]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[4]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[4]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[4]),
  .inena_out_mscbus(mp2_inena_out_mscbus[4]),
  .dir_out_mscbus(mp2_dir_out_mscbus[4]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[4]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[4]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[24:20]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[159:128]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[4]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[4]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[4]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[4]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[4]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[4]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[4]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[4]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[4]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_4_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_4_out_demux_peripheral_mscbus),
  .io_pad(MP2_4_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(289)) I_b_MP2_5(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[5]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[5]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[5]),
  .slew_out_mscbus(mp2_slew_out_mscbus[5]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[5]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[5]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[5]),
  .inena_out_mscbus(mp2_inena_out_mscbus[5]),
  .dir_out_mscbus(mp2_dir_out_mscbus[5]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[5]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[5]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[29:25]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[191:160]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[5]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[5]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[5]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[5]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[5]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[5]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[5]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[5]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[5]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_5_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_5_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP2_5_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(290)) I_b_MP2_6(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[6]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[6]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[6]),
  .slew_out_mscbus(mp2_slew_out_mscbus[6]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[6]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[6]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[6]),
  .inena_out_mscbus(mp2_inena_out_mscbus[6]),
  .dir_out_mscbus(mp2_dir_out_mscbus[6]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[6]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[6]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[34:30]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[223:192]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[6]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[6]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[6]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[6]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[6]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[6]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[6]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[6]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[6]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_6_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_6_out_demux_peripheral_mscbus),
  .io_pad(MP2_6_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(291)) I_b_MP2_7(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[7]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[7]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[7]),
  .slew_out_mscbus(mp2_slew_out_mscbus[7]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[7]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[7]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[7]),
  .inena_out_mscbus(mp2_inena_out_mscbus[7]),
  .dir_out_mscbus(mp2_dir_out_mscbus[7]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[7]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[7]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[39:35]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[255:224]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[7]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[7]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[7]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[7]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[7]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[7]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[7]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[7]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[7]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_7_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_7_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP2_7_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(292)) I_b_MP2_8(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[8]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[8]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[8]),
  .slew_out_mscbus(mp2_slew_out_mscbus[8]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[8]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[8]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[8]),
  .inena_out_mscbus(mp2_inena_out_mscbus[8]),
  .dir_out_mscbus(mp2_dir_out_mscbus[8]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[8]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[8]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[44:40]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[287:256]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[8]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[8]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[8]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[8]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[8]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[8]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[8]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[8]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[8]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_8_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_8_out_demux_peripheral_mscbus),
  .io_pad(MP2_8_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(293)) I_b_MP2_9(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[9]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[9]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[9]),
  .slew_out_mscbus(mp2_slew_out_mscbus[9]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[9]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[9]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[9]),
  .inena_out_mscbus(mp2_inena_out_mscbus[9]),
  .dir_out_mscbus(mp2_dir_out_mscbus[9]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[9]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[9]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[49:45]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[319:288]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[9]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[9]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[9]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[9]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[9]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[9]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[9]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[9]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[9]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP2_9_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP2_9_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP2_9_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(294)) I_b_MP2_10(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[10]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[10]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[10]),
  .slew_out_mscbus(mp2_slew_out_mscbus[10]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[10]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[10]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[10]),
  .inena_out_mscbus(mp2_inena_out_mscbus[10]),
  .dir_out_mscbus(mp2_dir_out_mscbus[10]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[10]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[10]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[54:50]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[351:320]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[10]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[10]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[10]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[10]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[10]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[10]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[10]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[10]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[10]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_10_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_10_out_demux_peripheral_mscbus),
  .io_pad(MP2_10_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(295)) I_b_MP2_11(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[11]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[11]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[11]),
  .slew_out_mscbus(mp2_slew_out_mscbus[11]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[11]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[11]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[11]),
  .inena_out_mscbus(mp2_inena_out_mscbus[11]),
  .dir_out_mscbus(mp2_dir_out_mscbus[11]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[11]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[11]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[59:55]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[383:352]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[11]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[11]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[11]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[11]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[11]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[11]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[11]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[11]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[11]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_11_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_11_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP2_11_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(2), .O_NUM_PERIPHERALS(2), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(296)) I_b_MP2_12(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[12]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[12]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[12]),
  .slew_out_mscbus(mp2_slew_out_mscbus[12]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[12]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[12]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[12]),
  .inena_out_mscbus(mp2_inena_out_mscbus[12]),
  .dir_out_mscbus(mp2_dir_out_mscbus[12]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[12]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[12]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[64:60]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[415:384]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[12]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[12]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[12]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[12]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[12]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[12]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[12]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[12]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[12]),
  .i_peripheral_oe({2{1'b1}}),
  .i_peripheral_out(MP2_12_in_mux_peripheral_mscbus[1:0]),
  .o_peripheral_in(MP2_12_out_demux_peripheral_mscbus[1:0]),
  .io_pad(MP2_12_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(297)) I_b_MP2_13(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[13]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[13]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[13]),
  .slew_out_mscbus(mp2_slew_out_mscbus[13]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[13]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[13]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[13]),
  .inena_out_mscbus(mp2_inena_out_mscbus[13]),
  .dir_out_mscbus(mp2_dir_out_mscbus[13]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[13]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[13]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[69:65]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[447:416]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[13]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[13]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[13]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[13]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[13]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[13]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[13]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[13]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[13]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP2_13_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP2_13_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP2_13_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(3), .O_NUM_PERIPHERALS(1), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(298)) I_b_MP2_14(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[14]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[14]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[14]),
  .slew_out_mscbus(mp2_slew_out_mscbus[14]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[14]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[14]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[14]),
  .inena_out_mscbus(mp2_inena_out_mscbus[14]),
  .dir_out_mscbus(mp2_dir_out_mscbus[14]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[14]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[14]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[74:70]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[479:448]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[14]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[14]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[14]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[14]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[14]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[14]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[14]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[14]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[14]),
  .i_peripheral_oe({3{1'b1}}),
  .i_peripheral_out(MP2_14_in_mux_peripheral_mscbus[2:0]),
  .o_peripheral_in(MP2_14_out_demux_peripheral_mscbus),
  .io_pad(MP2_14_IO)
);

pinmux_with_io_mp #(.I_NUM_PERIPHERALS(1), .O_NUM_PERIPHERALS(3), .DATA_WIDTH(1), .SEL_WIDTH(5), .array_cell_index(299)) I_b_MP2_15(
  .i_clk(gpio_clock),
  .i_clk_rc(clk_rc),
  .i_clk_perpll(clk_perpll),
  .i_rst_n(sys_reset_n),
  .amsel_out_mscbus(mp2_amsel_out_mscbus[15]),
  .ds0_out_mscbus(mp2_ds0_out_mscbus[15]),
  .ds1_out_mscbus(mp2_ds1_out_mscbus[15]),
  .slew_out_mscbus(mp2_slew_out_mscbus[15]),
  .schmitt_out_mscbus(mp2_schmitt_out_mscbus[15]),
  .mode0_out_mscbus(mp2_mode0_out_mscbus[15]),
  .mode1_out_mscbus(mp2_mode1_out_mscbus[15]),
  .inena_out_mscbus(mp2_inena_out_mscbus[15]),
  .dir_out_mscbus(mp2_dir_out_mscbus[15]),
  .pull_en_out_mscbus(mp2_pull_en_out_mscbus[15]),
  .pull_type_out_mscbus(mp2_pull_type_out_mscbus[15]),
  .pinmux_muxsel_out_mscbus(mp2_pinmux_muxsel_out_mscbus[79:75]),
  .in_function_en_out_mscbus(mp2_in_function_en_out_mscbus[511:480]),
  .async_in_from_pad_mscbus(mp2_async_in_from_pad_mscbus[15]),
  .gpio_out_2_buf_mscbus(mp2_gpio_out_2_buf_mscbus[15]),
  .gpio_out_en_2_buf_mscbus(mp2_gpio_out_en_2_buf_mscbus[15]),
  .pinmuxdata_2_gpio_mscbus(mp2_pinmuxdata_2_gpio_mscbus[15]),
  .pinmuxen_2_gpio_mscbus(mp2_pinmuxen_2_gpio_mscbus[15]),
  .GP_DATA_IN_out_mscbus(mp2_GP_DATA_IN_out_mscbus[15]),
  .data_out_2_pinmux_mscbus(mp2_data_out_2_pinmux_mscbus[15]),
  .lvds_en_ctrl_out_mscbus(mp2_lvds_en_ctrl_out_mscbus[15]),
  .in_termination_en_out_mscbus(mp2_in_termination_en_out_mscbus[15]),
  .i_peripheral_oe(1'b1),
  .i_peripheral_out(MP2_15_in_mux_peripheral_mscbus),
  .o_peripheral_in(MP2_15_out_demux_peripheral_mscbus[2:0]),
  .io_pad(MP2_15_IO)
);


endmodule


