//====================================================================
// Copyright (c) 2025 Texas Instruments, Inc.
// This is an unpublished work created in the year stated above.
// Texas Instruments owns all rights in and to this work and
// intends to maintain and protect it as an unpublished copyright.
// In the event of either inadvertent or deliberate publication,
// the above stated date shall be treated as the year of first
// publication. In the event of such publication, Texas Instruments
// intends to enforce its rights in the work under the copyright
// laws as a published work.
//====================================================================
//
// ioss_wrapper.v
//
//    ioss wrapper
//
//====================================================================
// Module Designer: Himanshi (h-himanshi@ti.com)
// Contact Info:    Texas Instruments
//                  DSP Systems /  Group
//                  12500 TI Blvd
//                  Dallas, Texas 75243
//                  (918)708-488241
//
//====================================================================
// Revision History:
//  1.0.0.0 15/1/2025 spec a0507242 first version
//
//====================================================================
// Generated by VeriPerl Compiler version 3.0.347
//    Build 2021.09.22.09.59.05
//
//====================================================================
`timescale 1 ps / 1 ps


module ioss_wrapper (

  // IO PORT
  AP0_IO,                                // I/O connection to toplevel

  // IO PORT
  AP1_IO,                                // I/O connection to toplevel

  // IO PORT
  AP10_IO,                               // I/O connection to toplevel

  // IO PORT
  AP11_IO,                               // I/O connection to toplevel

  // IO PORT
  AP12_IO,                               // I/O connection to toplevel

  // IO PORT
  AP13_IO,                               // I/O connection to toplevel

  // IO PORT
  AP14_IO,                               // I/O connection to toplevel

  // IO PORT
  AP15_IO,                               // I/O connection to toplevel

  // IO PORT
  AP16_IO,                               // I/O connection to toplevel

  // IO PORT
  AP17_IO,                               // I/O connection to toplevel

  // IO PORT
  AP18_IO,                               // I/O connection to toplevel

  // IO PORT
  AP19_IO,                               // I/O connection to toplevel

  // IO PORT
  AP2_IO,                                // I/O connection to toplevel

  // IO PORT
  AP20_IO,                               // I/O connection to toplevel

  // IO PORT
  AP21_IO,                               // I/O connection to toplevel

  // IO PORT
  AP22_IO,                               // I/O connection to toplevel

  // IO PORT
  AP23_IO,                               // I/O connection to toplevel

  // IO PORT
  AP24_IO,                               // I/O connection to toplevel

  // IO PORT
  AP25_IO,                               // I/O connection to toplevel

  // IO PORT
  AP26_IO,                               // I/O connection to toplevel

  // IO PORT
  AP27_IO,                               // I/O connection to toplevel

  // IO PORT
  AP28_IO,                               // I/O connection to toplevel

  // IO PORT
  AP29_IO,                               // I/O connection to toplevel

  // IO PORT
  AP3_IO,                                // I/O connection to toplevel

  // IO PORT
  AP30_IO,                               // I/O connection to toplevel

  // IO PORT
  AP31_IO,                               // I/O connection to toplevel

  // IO PORT
  AP32_IO,                               // I/O connection to toplevel

  // IO PORT
  AP33_IO,                               // I/O connection to toplevel

  // IO PORT
  AP34_IO,                               // I/O connection to toplevel

  // IO PORT
  AP35_IO,                               // I/O connection to toplevel

  // IO PORT
  AP36_IO,                               // I/O connection to toplevel

  // IO PORT
  AP37_IO,                               // I/O connection to toplevel

  // IO PORT
  AP38_IO,                               // I/O connection to toplevel

  // IO PORT
  AP39_IO,                               // I/O connection to toplevel

  // IO PORT
  AP4_IO,                                // I/O connection to toplevel

  // IO PORT
  AP40_IO,                               // I/O connection to toplevel

  // IO PORT
  AP41_IO,                               // I/O connection to toplevel

  // IO PORT
  AP42_IO,                               // I/O connection to toplevel

  // IO PORT
  AP43_IO,                               // I/O connection to toplevel

  // IO PORT
  AP44_IO,                               // I/O connection to toplevel

  // IO PORT
  AP45_IO,                               // I/O connection to toplevel

  // IO PORT
  AP46_IO,                               // I/O connection to toplevel

  // IO PORT
  AP47_IO,                               // I/O connection to toplevel

  // IO PORT
  AP5_IO,                                // I/O connection to toplevel

  // IO PORT
  AP6_IO,                                // I/O connection to toplevel

  // IO PORT
  AP7_IO,                                // I/O connection to toplevel

  // IO PORT
  AP8_IO,                                // I/O connection to toplevel

  // IO PORT
  AP9_IO,                                // I/O connection to toplevel

  // IO PORT
  AURORACLKN_IO,                         // I/O connection to toplevel

  // IO PORT
  AURORACLKP_IO,                         // I/O connection to toplevel

  // IO PORT
  AURORADN_IO,                           // I/O connection to toplevel

  // IO PORT
  AURORADP_IO,                           // I/O connection to toplevel

  // IO PORT
  DCDCNMOS_IO,                           // I/O connection to toplevel

  // IO PORT
  DCDCPMOS_IO,                           // I/O connection to toplevel

  // IO PORT
  DP0_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP0_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP0_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP1_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP1_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP2_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP2_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP3_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP3_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP4_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP4_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP5_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_28_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_29_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_30_IO,                             // I/O connection to toplevel

  // IO PORT
  DP5_31_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP6_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_15_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_16_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_17_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_18_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_19_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_20_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_21_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_22_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_23_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_24_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_25_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_26_IO,                             // I/O connection to toplevel

  // IO PORT
  DP6_27_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_0_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_1_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_2_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_3_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_4_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_5_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_6_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_7_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_8_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_9_IO,                              // I/O connection to toplevel

  // IO PORT
  DP7_10_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_11_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_12_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_13_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_14_IO,                             // I/O connection to toplevel

  // IO PORT
  DP7_15_IO,                             // I/O connection to toplevel

  // IO PORT
  ERROR_IO,                              // I/O connection to toplevel

  // IO PORT
  EXTPMICEN_IO,                          // I/O connection to toplevel

  // IO PORT
  FLASHTESTPAD1FT_IO,                    // I/O connection to toplevel

  // IO PORT
  FLASHTESTPAD2_IO,                      // I/O connection to toplevel

  // IO PORT
  FLASHTESTPAD3FT_IO,                    // I/O connection to toplevel

  // IO PORT
  FLASHTESTPAD4_IO,                      // I/O connection to toplevel

  // IO PORT
  FLASHTESTPAD5_IO,                      // I/O connection to toplevel

  // IO PORT
  MP0_0_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_1_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_2_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_3_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_4_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_5_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_6_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_7_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_8_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_9_IO,                              // I/O connection to toplevel

  // IO PORT
  MP0_10_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_11_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_12_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_13_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_14_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_15_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_16_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_17_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_18_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_19_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_20_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_21_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_22_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_23_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_24_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_25_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_26_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_27_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_28_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_29_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_30_IO,                             // I/O connection to toplevel

  // IO PORT
  MP0_31_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_0_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_1_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_2_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_3_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_4_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_5_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_6_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_7_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_8_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_9_IO,                              // I/O connection to toplevel

  // IO PORT
  MP1_10_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_11_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_12_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_13_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_14_IO,                             // I/O connection to toplevel

  // IO PORT
  MP1_15_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_0_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_1_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_2_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_3_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_4_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_5_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_6_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_7_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_8_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_9_IO,                              // I/O connection to toplevel

  // IO PORT
  MP2_10_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_11_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_12_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_13_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_14_IO,                             // I/O connection to toplevel

  // IO PORT
  MP2_15_IO,                             // I/O connection to toplevel

  // IO PORT
  PWR_ON_RSTn_IO,                        // I/O connection to toplevel

  // IO PORT
  RESETOUTn_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII0RXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII0RXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII0TXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII0TXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII1RXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII1RXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII1TXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII1TXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII2RXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII2RXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII2TXN_IO,                          // I/O connection to toplevel

  // IO PORT
  SGMII2TXP_IO,                          // I/O connection to toplevel

  // IO PORT
  SPI0LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI1LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI2LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI3LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI4LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI5LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI6LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI7LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI8LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  SPI9LPBCLKUNB_IO,                      // I/O connection to toplevel

  // IO PORT
  TCK_IO,                                // I/O connection to toplevel

  // IO PORT
  TDI_IO,                                // I/O connection to toplevel

  // IO PORT
  TDO_IO,                                // I/O connection to toplevel

  // IO PORT
  TMS_IO,                                // I/O connection to toplevel

  // IO PORT
  TRSTN_IO,                              // I/O connection to toplevel

  // IO PORT
  VDDS_REF_LPD_HI_IO,                    // I/O connection to toplevel

  // IO PORT
  VDDS_REF_LPD_LO_IO,                    // I/O connection to toplevel

  // IO PORT
  VDDS_REF_SD_HI_IO,                     // I/O connection to toplevel

  // IO PORT
  VDDS_REF_SD_LO_IO,                     // I/O connection to toplevel

  // IO PORT
  VDDS_REF0_HI_IO,                       // I/O connection to toplevel

  // IO PORT
  VDDS_REF0_LO_IO,                       // I/O connection to toplevel

  // IO PORT
  VDDS_REF1_HI_IO,                       // I/O connection to toplevel

  // IO PORT
  VDDS_REF1_LO_IO,                       // I/O connection to toplevel

  // IO PORT
  VDDS_REF2_HI_IO,                       // I/O connection to toplevel

  // IO PORT
  VDDS_REF2_LO_IO,                       // I/O connection to toplevel

  // IO PORT
  X1_IO,                                 // I/O connection to toplevel

  // IO PORT
  X2_IO,                                 // I/O connection to toplevel

  // IO PORT
  XSPI0LBCLKUNB_IO,                      // I/O connection to toplevel

  // PINMUX Clock interface
  pinmux_clock,                          // Module/peripheral clock

  // PINMUX Reset interface
  pinmux_reset_n,                        // Module/peripheral reset

  // GPIO Clock interface
  gpio_clock,                            // Module/peripheral clock

  // IO Clock interface
  io_clock,                              // Module/peripheral clock

  // IO Reset interface
  gpio_reset_n,                          // Module/peripheral reset

  // System Reset interface
  sys_reset_n,                           // Module/peripheral reset

  // IO Reset interface
  io_reset_n,                            // Module/peripheral reset

  // Clock Interface
  xbar_clk_clock,                        // Module/peripheral clock

  // Reset Interface
  xbar_rst_reset_n,                      // Module/peripheral reset

  // jtag_interface
  jtag_tck,                              // Clock
  jtag_trst_n,                           // Test reset
  jtag_tdi,                              // Data in
  jtag_tms,                              // State Select
  jtag_tdo_oe_n,                         // Data out enable
  jtag_tdo,                              // Data out

  // o_xrsn_pm_b_reset  interface
  o_xrsn_pm_b_reset_n,                   // Module/peripheral reset

  // o_xrsn_sw_fast_reset  interface
  o_xrsn_sw_fast_reset_n,                // Module/peripheral reset

  // o_porsn_frompmm_pm_d_reset  interface
  o_porsn_frompmm_pm_d_reset_n,          // Module/peripheral reset

  // o_porsn_pm_b_reset  interface
  o_porsn_pm_b_reset_n,                  // Module/peripheral reset

  // o_porsn_sw_pm_a_reset  interface
  o_porsn_sw_pm_a_reset_n,               // Module/peripheral reset

  // o_porsn_sw_pm_b_reset  interface
  o_porsn_sw_pm_b_reset_n,               // Module/peripheral reset

  // o_porsn_sw_pm_d_reset  interface
  o_porsn_sw_pm_d_reset_n,               // Module/peripheral reset

  // o_porsn_frompad_reset  interface
  o_porsn_frompad_reset_n,               // Module/peripheral reset

  // o_porsn_frompmm_pm_a_reset  interface
  o_porsn_frompmm_pm_a_reset_n,          // Module/peripheral reset

  // o_porsn_sw_streched_pm_a_reset  interface
  o_porsn_sw_streched_pm_a_reset_n,      // Module/peripheral reset

  // o_porsn_frompmm_pm_b_reset  interface
  o_porsn_frompmm_pm_b_reset_n,          // Module/peripheral reset

  // o_porsn_sw_streched_pm_b_reset  interface
  o_porsn_sw_streched_pm_b_reset_n,      // Module/peripheral reset

  // o_xrsn_frompad_reset  interface
  o_xrsn_frompad_reset_n,                // Module/peripheral reset

  // o_xrsn_sw_streched_reset  interface
  o_xrsn_sw_streched_reset_n,            // Module/peripheral reset

  // CBA_VBUSP_4_0 BUS Slave view interface
  io_vbusp_slv_routeid,                  // Route ID
  io_vbusp_slv_xid,                      // Transaction ID
  io_vbusp_slv_req,                      // Request
  io_vbusp_slv_dir,                      // Direction
  io_vbusp_slv_address,                  // Address
  io_vbusp_slv_xcnt,                     // Good Byte Count
  io_vbusp_slv_byten,                    // Byte Enables
  io_vbusp_slv_wdata,                    // Write Data
  io_vbusp_slv_wready,                   // Write Ready
  io_vbusp_slv_rdatap,                   // Read Data (Pipelined)
  io_vbusp_slv_rstatus,                  // Read Status
  io_vbusp_slv_rready,                   // Read Ready
  io_vbusp_slv_dtype,                    // Data Type
  io_vbusp_slv_priv,                     // Priviledge Attribute
  io_vbusp_slv_privid,                   // Priviledge ID
  io_vbusp_slv_secure,                   // Secure Attribute
  io_vbusp_slv_emudbg,                   // Emulation Debug Attribute

  // LPD_CAN0TX interface
  io_LPD_CAN0TX_txd,                     // CAN bus Transmit Data
  io_LPD_CAN0TX_rxd,                     // CAN bus Receive Data

  // LPD_CAN0RX interface
  io_LPD_CAN0RX_txd,                     // CAN bus Transmit Data
  io_LPD_CAN0RX_rxd,                     // CAN bus Receive Data

  // LPD_LIN0TX interface
  io_LPD_LIN0TX_txd,                     // Serial Data Transmission
  io_LPD_LIN0TX_rxd,                     // Serial Data Reception
  io_LPD_LIN0TX_tr_en,                   // Transceiver enable

  // LPD_LIN0RX interface
  io_LPD_LIN0RX_txd,                     // Serial Data Transmission
  io_LPD_LIN0RX_rxd,                     // Serial Data Reception
  io_LPD_LIN0RX_tr_en,                   // Transceiver enable

  // EPWM0 interface
  io_EPWM0_a_i,                          
  io_EPWM0_a_o,                          
  io_EPWM0_a_oen,                        
  io_EPWM0_b_i,                          
  io_EPWM0_b_o,                          
  io_EPWM0_b_oen,                        

  // EPWM1 interface
  io_EPWM1_a_i,                          
  io_EPWM1_a_o,                          
  io_EPWM1_a_oen,                        
  io_EPWM1_b_i,                          
  io_EPWM1_b_o,                          
  io_EPWM1_b_oen,                        

  // EPWM2 interface
  io_EPWM2_a_i,                          
  io_EPWM2_a_o,                          
  io_EPWM2_a_oen,                        
  io_EPWM2_b_i,                          
  io_EPWM2_b_o,                          
  io_EPWM2_b_oen,                        

  // EPWM3 interface
  io_EPWM3_a_i,                          
  io_EPWM3_a_o,                          
  io_EPWM3_a_oen,                        
  io_EPWM3_b_i,                          
  io_EPWM3_b_o,                          
  io_EPWM3_b_oen,                        

  // EPWM4 interface
  io_EPWM4_a_i,                          
  io_EPWM4_a_o,                          
  io_EPWM4_a_oen,                        
  io_EPWM4_b_i,                          
  io_EPWM4_b_o,                          
  io_EPWM4_b_oen,                        

  // EPWM5 interface
  io_EPWM5_a_i,                          
  io_EPWM5_a_o,                          
  io_EPWM5_a_oen,                        
  io_EPWM5_b_i,                          
  io_EPWM5_b_o,                          
  io_EPWM5_b_oen,                        

  // EPWM6 interface
  io_EPWM6_a_i,                          
  io_EPWM6_a_o,                          
  io_EPWM6_a_oen,                        
  io_EPWM6_b_i,                          
  io_EPWM6_b_o,                          
  io_EPWM6_b_oen,                        

  // EPWM7 interface
  io_EPWM7_a_i,                          
  io_EPWM7_a_o,                          
  io_EPWM7_a_oen,                        
  io_EPWM7_b_i,                          
  io_EPWM7_b_o,                          
  io_EPWM7_b_oen,                        

  // EPWM8 interface
  io_EPWM8_a_i,                          
  io_EPWM8_a_o,                          
  io_EPWM8_a_oen,                        
  io_EPWM8_b_i,                          
  io_EPWM8_b_o,                          
  io_EPWM8_b_oen,                        

  // EPWM9 interface
  io_EPWM9_a_i,                          
  io_EPWM9_a_o,                          
  io_EPWM9_a_oen,                        
  io_EPWM9_b_i,                          
  io_EPWM9_b_o,                          
  io_EPWM9_b_oen,                        

  // EPWM10 interface
  io_EPWM10_a_i,                         
  io_EPWM10_a_o,                         
  io_EPWM10_a_oen,                       
  io_EPWM10_b_i,                         
  io_EPWM10_b_o,                         
  io_EPWM10_b_oen,                       

  // EPWM11 interface
  io_EPWM11_a_i,                         
  io_EPWM11_a_o,                         
  io_EPWM11_a_oen,                       
  io_EPWM11_b_i,                         
  io_EPWM11_b_o,                         
  io_EPWM11_b_oen,                       

  // EPWM12 interface
  io_EPWM12_a_i,                         
  io_EPWM12_a_o,                         
  io_EPWM12_a_oen,                       
  io_EPWM12_b_i,                         
  io_EPWM12_b_o,                         
  io_EPWM12_b_oen,                       

  // EPWM13 interface
  io_EPWM13_a_i,                         
  io_EPWM13_a_o,                         
  io_EPWM13_a_oen,                       
  io_EPWM13_b_i,                         
  io_EPWM13_b_o,                         
  io_EPWM13_b_oen,                       

  // EPWM14 interface
  io_EPWM14_a_i,                         
  io_EPWM14_a_o,                         
  io_EPWM14_a_oen,                       
  io_EPWM14_b_i,                         
  io_EPWM14_b_o,                         
  io_EPWM14_b_oen,                       

  // EPWM15 interface
  io_EPWM15_a_i,                         
  io_EPWM15_a_o,                         
  io_EPWM15_a_oen,                       
  io_EPWM15_b_i,                         
  io_EPWM15_b_o,                         
  io_EPWM15_b_oen,                       

  // EPWM16 interface
  io_EPWM16_a_i,                         
  io_EPWM16_a_o,                         
  io_EPWM16_a_oen,                       
  io_EPWM16_b_i,                         
  io_EPWM16_b_o,                         
  io_EPWM16_b_oen,                       

  // EPWM17 interface
  io_EPWM17_a_i,                         
  io_EPWM17_a_o,                         
  io_EPWM17_a_oen,                       
  io_EPWM17_b_i,                         
  io_EPWM17_b_o,                         
  io_EPWM17_b_oen,                       

  // EPWM18 interface
  io_EPWM18_a_i,                         
  io_EPWM18_a_o,                         
  io_EPWM18_a_oen,                       
  io_EPWM18_b_i,                         
  io_EPWM18_b_o,                         
  io_EPWM18_b_oen,                       

  // EPWM19 interface
  io_EPWM19_a_i,                         
  io_EPWM19_a_o,                         
  io_EPWM19_a_oen,                       
  io_EPWM19_b_i,                         
  io_EPWM19_b_o,                         
  io_EPWM19_b_oen,                       

  // EPWM20 interface
  io_EPWM20_a_i,                         
  io_EPWM20_a_o,                         
  io_EPWM20_a_oen,                       
  io_EPWM20_b_i,                         
  io_EPWM20_b_o,                         
  io_EPWM20_b_oen,                       

  // EPWM21 interface
  io_EPWM21_a_i,                         
  io_EPWM21_a_o,                         
  io_EPWM21_a_oen,                       
  io_EPWM21_b_i,                         
  io_EPWM21_b_o,                         
  io_EPWM21_b_oen,                       

  // EPWM22 interface
  io_EPWM22_a_i,                         
  io_EPWM22_a_o,                         
  io_EPWM22_a_oen,                       
  io_EPWM22_b_i,                         
  io_EPWM22_b_o,                         
  io_EPWM22_b_oen,                       

  // EPWM23 interface
  io_EPWM23_a_i,                         
  io_EPWM23_a_o,                         
  io_EPWM23_a_oen,                       
  io_EPWM23_b_i,                         
  io_EPWM23_b_o,                         
  io_EPWM23_b_oen,                       

  // EPWM24 interface
  io_EPWM24_a_i,                         
  io_EPWM24_a_o,                         
  io_EPWM24_a_oen,                       
  io_EPWM24_b_i,                         
  io_EPWM24_b_o,                         
  io_EPWM24_b_oen,                       

  // EPWM25 interface
  io_EPWM25_a_i,                         
  io_EPWM25_a_o,                         
  io_EPWM25_a_oen,                       
  io_EPWM25_b_i,                         
  io_EPWM25_b_o,                         
  io_EPWM25_b_oen,                       

  // EPWM26 interface
  io_EPWM26_a_i,                         
  io_EPWM26_a_o,                         
  io_EPWM26_a_oen,                       
  io_EPWM26_b_i,                         
  io_EPWM26_b_o,                         
  io_EPWM26_b_oen,                       

  // EPWM27 interface
  io_EPWM27_a_i,                         
  io_EPWM27_a_o,                         
  io_EPWM27_a_oen,                       
  io_EPWM27_b_i,                         
  io_EPWM27_b_o,                         
  io_EPWM27_b_oen,                       

  // EPWM28 interface
  io_EPWM28_a_i,                         
  io_EPWM28_a_o,                         
  io_EPWM28_a_oen,                       
  io_EPWM28_b_i,                         
  io_EPWM28_b_o,                         
  io_EPWM28_b_oen,                       

  // EPWM29 interface
  io_EPWM29_a_i,                         
  io_EPWM29_a_o,                         
  io_EPWM29_a_oen,                       
  io_EPWM29_b_i,                         
  io_EPWM29_b_o,                         
  io_EPWM29_b_oen,                       

  // EPWM30 interface
  io_EPWM30_a_i,                         
  io_EPWM30_a_o,                         
  io_EPWM30_a_oen,                       
  io_EPWM30_b_i,                         
  io_EPWM30_b_o,                         
  io_EPWM30_b_oen,                       

  // EPWM31 interface
  io_EPWM31_a_i,                         
  io_EPWM31_a_o,                         
  io_EPWM31_a_oen,                       
  io_EPWM31_b_i,                         
  io_EPWM31_b_o,                         
  io_EPWM31_b_oen,                       

  // EPWMSYNCO interface
  io_EPWMSYNCO_a_i,                      
  io_EPWMSYNCO_a_o,                      
  io_EPWMSYNCO_a_oen,                    
  io_EPWMSYNCO_b_i,                      
  io_EPWMSYNCO_b_o,                      
  io_EPWMSYNCO_b_oen,                    

  // ICL  PORT
  io_OUTPUTXBAR0_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR1_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR2_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR3_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR4_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR5_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR6_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR7_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR8_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR9_intr,                   // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR10_intr,                  // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR11_intr,                  // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR12_intr,                  // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR13_intr,                  // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR14_intr,                  // Interrupt signal

  // ICL  PORT
  io_OUTPUTXBAR15_intr,                  // Interrupt signal

  // SDFM_SDFM0 interface
  io_SDFM0_i_datain1,                    // DATAIN1
  io_SDFM0_i_clock1,                     // CLOCK1
  io_SDFM0_i_datain2,                    // DATAIN2
  io_SDFM0_i_clock2,                     // CLOCK2
  io_SDFM0_i_datain3,                    // DATAIN3
  io_SDFM0_i_clock3,                     // CLOCK3
  io_SDFM0_i_datain4,                    // DATAIN4
  io_SDFM0_i_clock4,                     // CLOCK4

  // SDFM_SDFM1 interface
  io_SDFM1_i_datain1,                    // DATAIN1
  io_SDFM1_i_clock1,                     // CLOCK1
  io_SDFM1_i_datain2,                    // DATAIN2
  io_SDFM1_i_clock2,                     // CLOCK2
  io_SDFM1_i_datain3,                    // DATAIN3
  io_SDFM1_i_clock3,                     // CLOCK3
  io_SDFM1_i_datain4,                    // DATAIN4
  io_SDFM1_i_clock4,                     // CLOCK4

  // SDFM_SDFM2 interface
  io_SDFM2_i_datain1,                    // DATAIN1
  io_SDFM2_i_clock1,                     // CLOCK1
  io_SDFM2_i_datain2,                    // DATAIN2
  io_SDFM2_i_clock2,                     // CLOCK2
  io_SDFM2_i_datain3,                    // DATAIN3
  io_SDFM2_i_clock3,                     // CLOCK3
  io_SDFM2_i_datain4,                    // DATAIN4
  io_SDFM2_i_clock4,                     // CLOCK4

  // SDFM_SDFM3 interface
  io_SDFM3_i_datain1,                    // DATAIN1
  io_SDFM3_i_clock1,                     // CLOCK1
  io_SDFM3_i_datain2,                    // DATAIN2
  io_SDFM3_i_clock2,                     // CLOCK2
  io_SDFM3_i_datain3,                    // DATAIN3
  io_SDFM3_i_clock3,                     // CLOCK3
  io_SDFM3_i_datain4,                    // DATAIN4
  io_SDFM3_i_clock4,                     // CLOCK4

  // SDFM_SDFM4 interface
  io_SDFM4_i_datain1,                    // DATAIN1
  io_SDFM4_i_clock1,                     // CLOCK1
  io_SDFM4_i_datain2,                    // DATAIN2
  io_SDFM4_i_clock2,                     // CLOCK2
  io_SDFM4_i_datain3,                    // DATAIN3
  io_SDFM4_i_clock3,                     // CLOCK3
  io_SDFM4_i_datain4,                    // DATAIN4
  io_SDFM4_i_clock4,                     // CLOCK4

  // SDFM_SDFM5 interface
  io_SDFM5_i_datain1,                    // DATAIN1
  io_SDFM5_i_clock1,                     // CLOCK1
  io_SDFM5_i_datain2,                    // DATAIN2
  io_SDFM5_i_clock2,                     // CLOCK2
  io_SDFM5_i_datain3,                    // DATAIN3
  io_SDFM5_i_clock3,                     // CLOCK3
  io_SDFM5_i_datain4,                    // DATAIN4
  io_SDFM5_i_clock4,                     // CLOCK4

  // SDFM_SDFM6 interface
  io_SDFM6_i_datain1,                    // DATAIN1
  io_SDFM6_i_clock1,                     // CLOCK1
  io_SDFM6_i_datain2,                    // DATAIN2
  io_SDFM6_i_clock2,                     // CLOCK2
  io_SDFM6_i_datain3,                    // DATAIN3
  io_SDFM6_i_clock3,                     // CLOCK3
  io_SDFM6_i_datain4,                    // DATAIN4
  io_SDFM6_i_clock4,                     // CLOCK4

  // SDFM_SDFM7 interface
  io_SDFM7_i_datain1,                    // DATAIN1
  io_SDFM7_i_clock1,                     // CLOCK1
  io_SDFM7_i_datain2,                    // DATAIN2
  io_SDFM7_i_clock2,                     // CLOCK2
  io_SDFM7_i_datain3,                    // DATAIN3
  io_SDFM7_i_clock3,                     // CLOCK3
  io_SDFM7_i_datain4,                    // DATAIN4
  io_SDFM7_i_clock4,                     // CLOCK4

  // SDFM_SDFM8 interface
  io_SDFM8_i_datain1,                    // DATAIN1
  io_SDFM8_i_clock1,                     // CLOCK1
  io_SDFM8_i_datain2,                    // DATAIN2
  io_SDFM8_i_clock2,                     // CLOCK2
  io_SDFM8_i_datain3,                    // DATAIN3
  io_SDFM8_i_clock3,                     // CLOCK3
  io_SDFM8_i_datain4,                    // DATAIN4
  io_SDFM8_i_clock4,                     // CLOCK4

  // SDFM_SDFM9 interface
  io_SDFM9_i_datain1,                    // DATAIN1
  io_SDFM9_i_clock1,                     // CLOCK1
  io_SDFM9_i_datain2,                    // DATAIN2
  io_SDFM9_i_clock2,                     // CLOCK2
  io_SDFM9_i_datain3,                    // DATAIN3
  io_SDFM9_i_clock3,                     // CLOCK3
  io_SDFM9_i_datain4,                    // DATAIN4
  io_SDFM9_i_clock4,                     // CLOCK4

  // SDFM_SDFM10 interface
  io_SDFM10_i_datain1,                   // DATAIN1
  io_SDFM10_i_clock1,                    // CLOCK1
  io_SDFM10_i_datain2,                   // DATAIN2
  io_SDFM10_i_clock2,                    // CLOCK2
  io_SDFM10_i_datain3,                   // DATAIN3
  io_SDFM10_i_clock3,                    // CLOCK3
  io_SDFM10_i_datain4,                   // DATAIN4
  io_SDFM10_i_clock4,                    // CLOCK4

  // SDFM_SDFM11 interface
  io_SDFM11_i_datain1,                   // DATAIN1
  io_SDFM11_i_clock1,                    // CLOCK1
  io_SDFM11_i_datain2,                   // DATAIN2
  io_SDFM11_i_clock2,                    // CLOCK2
  io_SDFM11_i_datain3,                   // DATAIN3
  io_SDFM11_i_clock3,                    // CLOCK3
  io_SDFM11_i_datain4,                   // DATAIN4
  io_SDFM11_i_clock4,                    // CLOCK4

  // ADC0EXTMUXSEL0 interface
  io_ADC0EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC0EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC0EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC0EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC0EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC0EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC0EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC0EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC0EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC0EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC0EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC0EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC0EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC0EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC0EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC0EXTMUXSEL0 interface
  io_ext_ADC0EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC0EXTMUXSEL1 interface
  io_ADC0EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC0EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC0EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC0EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC0EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC0EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC0EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC0EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC0EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC0EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC0EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC0EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC0EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC0EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC0EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC0EXTMUXSEL1 interface
  io_ext_ADC0EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC0EXTMUXSEL2 interface
  io_ADC0EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC0EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC0EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC0EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC0EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC0EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC0EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC0EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC0EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC0EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC0EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC0EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC0EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC0EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC0EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC0EXTMUXSEL2 interface
  io_ext_ADC0EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC0EXTMUXSEL3 interface
  io_ADC0EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC0EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC0EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC0EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC0EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC0EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC0EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC0EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC0EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC0EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC0EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC0EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC0EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC0EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC0EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC0EXTMUXSEL3 interface
  io_ext_ADC0EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC1EXTMUXSEL0 interface
  io_ADC1EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC1EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC1EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC1EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC1EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC1EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC1EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC1EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC1EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC1EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC1EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC1EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC1EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC1EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC1EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC1EXTMUXSEL0 interface
  io_ext_ADC1EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC1EXTMUXSEL1 interface
  io_ADC1EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC1EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC1EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC1EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC1EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC1EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC1EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC1EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC1EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC1EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC1EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC1EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC1EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC1EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC1EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC1EXTMUXSEL1 interface
  io_ext_ADC1EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC1EXTMUXSEL2 interface
  io_ADC1EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC1EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC1EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC1EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC1EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC1EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC1EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC1EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC1EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC1EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC1EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC1EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC1EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC1EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC1EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC1EXTMUXSEL2 interface
  io_ext_ADC1EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC1EXTMUXSEL3 interface
  io_ADC1EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC1EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC1EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC1EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC1EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC1EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC1EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC1EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC1EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC1EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC1EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC1EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC1EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC1EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC1EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC1EXTMUXSEL3 interface
  io_ext_ADC1EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC2EXTMUXSEL0 interface
  io_ADC2EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC2EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC2EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC2EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC2EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC2EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC2EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC2EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC2EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC2EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC2EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC2EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC2EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC2EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC2EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC2EXTMUXSEL0 interface
  io_ext_ADC2EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC2EXTMUXSEL1 interface
  io_ADC2EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC2EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC2EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC2EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC2EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC2EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC2EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC2EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC2EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC2EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC2EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC2EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC2EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC2EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC2EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC2EXTMUXSEL1 interface
  io_ext_ADC2EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC2EXTMUXSEL2 interface
  io_ADC2EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC2EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC2EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC2EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC2EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC2EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC2EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC2EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC2EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC2EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC2EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC2EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC2EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC2EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC2EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC2EXTMUXSEL2 interface
  io_ext_ADC2EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC2EXTMUXSEL3 interface
  io_ADC2EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC2EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC2EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC2EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC2EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC2EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC2EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC2EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC2EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC2EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC2EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC2EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC2EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC2EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC2EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC2EXTMUXSEL3 interface
  io_ext_ADC2EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC3EXTMUXSEL0 interface
  io_ADC3EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC3EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC3EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC3EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC3EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC3EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC3EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC3EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC3EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC3EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC3EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC3EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC3EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC3EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC3EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC3EXTMUXSEL0 interface
  io_ext_ADC3EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC3EXTMUXSEL1 interface
  io_ADC3EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC3EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC3EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC3EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC3EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC3EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC3EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC3EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC3EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC3EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC3EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC3EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC3EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC3EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC3EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC3EXTMUXSEL1 interface
  io_ext_ADC3EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC3EXTMUXSEL2 interface
  io_ADC3EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC3EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC3EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC3EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC3EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC3EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC3EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC3EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC3EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC3EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC3EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC3EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC3EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC3EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC3EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC3EXTMUXSEL2 interface
  io_ext_ADC3EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC3EXTMUXSEL3 interface
  io_ADC3EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC3EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC3EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC3EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC3EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC3EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC3EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC3EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC3EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC3EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC3EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC3EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC3EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC3EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC3EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC3EXTMUXSEL3 interface
  io_ext_ADC3EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC4EXTMUXSEL0 interface
  io_ADC4EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC4EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC4EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC4EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC4EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC4EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC4EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC4EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC4EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC4EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC4EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC4EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC4EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC4EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC4EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC4EXTMUXSEL0 interface
  io_ext_ADC4EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC4EXTMUXSEL1 interface
  io_ADC4EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC4EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC4EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC4EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC4EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC4EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC4EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC4EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC4EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC4EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC4EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC4EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC4EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC4EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC4EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC4EXTMUXSEL1 interface
  io_ext_ADC4EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC4EXTMUXSEL2 interface
  io_ADC4EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC4EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC4EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC4EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC4EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC4EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC4EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC4EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC4EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC4EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC4EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC4EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC4EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC4EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC4EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC4EXTMUXSEL2 interface
  io_ext_ADC4EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC4EXTMUXSEL3 interface
  io_ADC4EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC4EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC4EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC4EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC4EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC4EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC4EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC4EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC4EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC4EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC4EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC4EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC4EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC4EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC4EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC4EXTMUXSEL3 interface
  io_ext_ADC4EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC5EXTMUXSEL0 interface
  io_ADC5EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC5EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC5EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC5EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC5EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC5EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC5EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC5EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC5EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC5EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC5EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC5EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC5EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC5EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC5EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC5EXTMUXSEL0 interface
  io_ext_ADC5EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC5EXTMUXSEL1 interface
  io_ADC5EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC5EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC5EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC5EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC5EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC5EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC5EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC5EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC5EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC5EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC5EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC5EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC5EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC5EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC5EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC5EXTMUXSEL1 interface
  io_ext_ADC5EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC5EXTMUXSEL2 interface
  io_ADC5EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC5EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC5EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC5EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC5EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC5EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC5EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC5EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC5EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC5EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC5EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC5EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC5EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC5EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC5EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC5EXTMUXSEL2 interface
  io_ext_ADC5EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC5EXTMUXSEL3 interface
  io_ADC5EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC5EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC5EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC5EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC5EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC5EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC5EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC5EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC5EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC5EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC5EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC5EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC5EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC5EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC5EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC5EXTMUXSEL3 interface
  io_ext_ADC5EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC6EXTMUXSEL0 interface
  io_ADC6EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC6EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC6EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC6EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC6EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC6EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC6EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC6EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC6EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC6EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC6EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC6EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC6EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC6EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC6EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC6EXTMUXSEL0 interface
  io_ext_ADC6EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC6EXTMUXSEL1 interface
  io_ADC6EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC6EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC6EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC6EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC6EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC6EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC6EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC6EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC6EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC6EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC6EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC6EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC6EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC6EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC6EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC6EXTMUXSEL1 interface
  io_ext_ADC6EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC6EXTMUXSEL2 interface
  io_ADC6EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC6EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC6EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC6EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC6EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC6EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC6EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC6EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC6EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC6EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC6EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC6EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC6EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC6EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC6EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC6EXTMUXSEL2 interface
  io_ext_ADC6EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC6EXTMUXSEL3 interface
  io_ADC6EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC6EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC6EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC6EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC6EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC6EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC6EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC6EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC6EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC6EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC6EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC6EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC6EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC6EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC6EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC6EXTMUXSEL3 interface
  io_ext_ADC6EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADC7EXTMUXSEL0 interface
  io_ADC7EXTMUXSEL0_adcconfig,           // ADC Config to ADC
  io_ADC7EXTMUXSEL0_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC7EXTMUXSEL0_adcofftrim,          // ADC Offset trim to ADC
  io_ADC7EXTMUXSEL0_adcresult,           // 16 bit result from ADC
  io_ADC7EXTMUXSEL0_adcclk,              // Divided clock to ADC.
  io_ADC7EXTMUXSEL0_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC7EXTMUXSEL0_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC7EXTMUXSEL0_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC7EXTMUXSEL0_adcpwrdn,            // ADC power down signal.
  io_ADC7EXTMUXSEL0_adcchsel,            // ADC Channel number to be converted.
  io_ADC7EXTMUXSEL0_adccalibmode,        // ADC calibmode
  io_ADC7EXTMUXSEL0_adccalibstep,        // ADC calibstep
  io_ADC7EXTMUXSEL0_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC7EXTMUXSEL0_samcapreset_level,   // ADC Sampcapreset level
  io_ADC7EXTMUXSEL0_dtb,                 // DTB bits for debug

  // ext_ADC7EXTMUXSEL0 interface
  io_ext_ADC7EXTMUXSEL0_adcchsel,        // ADC Channel number to be converted.

  // ADC7EXTMUXSEL1 interface
  io_ADC7EXTMUXSEL1_adcconfig,           // ADC Config to ADC
  io_ADC7EXTMUXSEL1_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC7EXTMUXSEL1_adcofftrim,          // ADC Offset trim to ADC
  io_ADC7EXTMUXSEL1_adcresult,           // 16 bit result from ADC
  io_ADC7EXTMUXSEL1_adcclk,              // Divided clock to ADC.
  io_ADC7EXTMUXSEL1_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC7EXTMUXSEL1_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC7EXTMUXSEL1_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC7EXTMUXSEL1_adcpwrdn,            // ADC power down signal.
  io_ADC7EXTMUXSEL1_adcchsel,            // ADC Channel number to be converted.
  io_ADC7EXTMUXSEL1_adccalibmode,        // ADC calibmode
  io_ADC7EXTMUXSEL1_adccalibstep,        // ADC calibstep
  io_ADC7EXTMUXSEL1_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC7EXTMUXSEL1_samcapreset_level,   // ADC Sampcapreset level
  io_ADC7EXTMUXSEL1_dtb,                 // DTB bits for debug

  // ext_ADC7EXTMUXSEL1 interface
  io_ext_ADC7EXTMUXSEL1_adcchsel,        // ADC Channel number to be converted.

  // ADC7EXTMUXSEL2 interface
  io_ADC7EXTMUXSEL2_adcconfig,           // ADC Config to ADC
  io_ADC7EXTMUXSEL2_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC7EXTMUXSEL2_adcofftrim,          // ADC Offset trim to ADC
  io_ADC7EXTMUXSEL2_adcresult,           // 16 bit result from ADC
  io_ADC7EXTMUXSEL2_adcclk,              // Divided clock to ADC.
  io_ADC7EXTMUXSEL2_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC7EXTMUXSEL2_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC7EXTMUXSEL2_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC7EXTMUXSEL2_adcpwrdn,            // ADC power down signal.
  io_ADC7EXTMUXSEL2_adcchsel,            // ADC Channel number to be converted.
  io_ADC7EXTMUXSEL2_adccalibmode,        // ADC calibmode
  io_ADC7EXTMUXSEL2_adccalibstep,        // ADC calibstep
  io_ADC7EXTMUXSEL2_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC7EXTMUXSEL2_samcapreset_level,   // ADC Sampcapreset level
  io_ADC7EXTMUXSEL2_dtb,                 // DTB bits for debug

  // ext_ADC7EXTMUXSEL2 interface
  io_ext_ADC7EXTMUXSEL2_adcchsel,        // ADC Channel number to be converted.

  // ADC7EXTMUXSEL3 interface
  io_ADC7EXTMUXSEL3_adcconfig,           // ADC Config to ADC
  io_ADC7EXTMUXSEL3_adcinltrim1,         // ADC Linearity Trim 1 to ADC
  io_ADC7EXTMUXSEL3_adcofftrim,          // ADC Offset trim to ADC
  io_ADC7EXTMUXSEL3_adcresult,           // 16 bit result from ADC
  io_ADC7EXTMUXSEL3_adcclk,              // Divided clock to ADC.
  io_ADC7EXTMUXSEL3_adcresolution,       // 16 bit / 12 bit resolution
  io_ADC7EXTMUXSEL3_adcsignalmode,       // Single ended Vs Differential mode
  io_ADC7EXTMUXSEL3_adcsoc,              // ADC start of conversion signal to ADC.
  io_ADC7EXTMUXSEL3_adcpwrdn,            // ADC power down signal.
  io_ADC7EXTMUXSEL3_adcchsel,            // ADC Channel number to be converted.
  io_ADC7EXTMUXSEL3_adccalibmode,        // ADC calibmode
  io_ADC7EXTMUXSEL3_adccalibstep,        // ADC calibstep
  io_ADC7EXTMUXSEL3_samcapreset_disable, // ADC Sampcapreset disable
  io_ADC7EXTMUXSEL3_samcapreset_level,   // ADC Sampcapreset level
  io_ADC7EXTMUXSEL3_dtb,                 // DTB bits for debug

  // ext_ADC7EXTMUXSEL3 interface
  io_ext_ADC7EXTMUXSEL3_adcchsel,        // ADC Channel number to be converted.

  // ADCSOC0 interface
  io_ADCSOC0_adcconfig,                  // ADC Config to ADC
  io_ADCSOC0_adcinltrim1,                // ADC Linearity Trim 1 to ADC
  io_ADCSOC0_adcofftrim,                 // ADC Offset trim to ADC
  io_ADCSOC0_adcresult,                  // 16 bit result from ADC
  io_ADCSOC0_adcclk,                     // Divided clock to ADC.
  io_ADCSOC0_adcresolution,              // 16 bit / 12 bit resolution
  io_ADCSOC0_adcsignalmode,              // Single ended Vs Differential mode
  io_ADCSOC0_adcsoc,                     // ADC start of conversion signal to ADC.
  io_ADCSOC0_adcpwrdn,                   // ADC power down signal.
  io_ADCSOC0_adcchsel,                   // ADC Channel number to be converted.
  io_ADCSOC0_adccalibmode,               // ADC calibmode
  io_ADCSOC0_adccalibstep,               // ADC calibstep
  io_ADCSOC0_samcapreset_disable,        // ADC Sampcapreset disable
  io_ADCSOC0_samcapreset_level,          // ADC Sampcapreset level
  io_ADCSOC0_dtb,                        // DTB bits for debug

  // ext_ADCSOC0 interface
  io_ext_ADCSOC0_adcchsel,               // ADC Channel number to be converted.

  // ADCSOC1 interface
  io_ADCSOC1_adcconfig,                  // ADC Config to ADC
  io_ADCSOC1_adcinltrim1,                // ADC Linearity Trim 1 to ADC
  io_ADCSOC1_adcofftrim,                 // ADC Offset trim to ADC
  io_ADCSOC1_adcresult,                  // 16 bit result from ADC
  io_ADCSOC1_adcclk,                     // Divided clock to ADC.
  io_ADCSOC1_adcresolution,              // 16 bit / 12 bit resolution
  io_ADCSOC1_adcsignalmode,              // Single ended Vs Differential mode
  io_ADCSOC1_adcsoc,                     // ADC start of conversion signal to ADC.
  io_ADCSOC1_adcpwrdn,                   // ADC power down signal.
  io_ADCSOC1_adcchsel,                   // ADC Channel number to be converted.
  io_ADCSOC1_adccalibmode,               // ADC calibmode
  io_ADCSOC1_adccalibstep,               // ADC calibstep
  io_ADCSOC1_samcapreset_disable,        // ADC Sampcapreset disable
  io_ADCSOC1_samcapreset_level,          // ADC Sampcapreset level
  io_ADCSOC1_dtb,                        // DTB bits for debug

  // ext_ADCSOC1 interface
  io_ext_ADCSOC1_adcchsel,               // ADC Channel number to be converted.

  // FSI0TX interface
  io_FSI0TX_ck,                          // Clock
  io_FSI0TX_d0,                          // Data0
  io_FSI0TX_d1,                          // Data1

  // FSI0RX interface
  io_FSI0RX_ck,                          // Clock
  io_FSI0RX_d0,                          // Data0
  io_FSI0RX_d1,                          // Data1

  // FSI1TX interface
  io_FSI1TX_ck,                          // Clock
  io_FSI1TX_d0,                          // Data0
  io_FSI1TX_d1,                          // Data1

  // FSI1RX interface
  io_FSI1RX_ck,                          // Clock
  io_FSI1RX_d0,                          // Data0
  io_FSI1RX_d1,                          // Data1

  // FSI2TX interface
  io_FSI2TX_ck,                          // Clock
  io_FSI2TX_d0,                          // Data0
  io_FSI2TX_d1,                          // Data1

  // FSI2RX interface
  io_FSI2RX_ck,                          // Clock
  io_FSI2RX_d0,                          // Data0
  io_FSI2RX_d1,                          // Data1

  // FSI3TX interface
  io_FSI3TX_ck,                          // Clock
  io_FSI3TX_d0,                          // Data0
  io_FSI3TX_d1,                          // Data1

  // FSI3RX interface
  io_FSI3RX_ck,                          // Clock
  io_FSI3RX_d0,                          // Data0
  io_FSI3RX_d1,                          // Data1

  // FSI4TX interface
  io_FSI4TX_ck,                          // Clock
  io_FSI4TX_d0,                          // Data0
  io_FSI4TX_d1,                          // Data1

  // FSI4RX interface
  io_FSI4RX_ck,                          // Clock
  io_FSI4RX_d0,                          // Data0
  io_FSI4RX_d1,                          // Data1

  // FSI5TX interface
  io_FSI5TX_ck,                          // Clock
  io_FSI5TX_d0,                          // Data0
  io_FSI5TX_d1,                          // Data1

  // FSI5RX interface
  io_FSI5RX_ck,                          // Clock
  io_FSI5RX_d0,                          // Data0
  io_FSI5RX_d1,                          // Data1

  // I2C0SCL interface
  io_I2C0SCL_piscl,                      // SCL input
  io_I2C0SCL_pisda,                      // SDA input
  io_I2C0SCL_porscl,                     // SCL output
  io_I2C0SCL_porsda,                     // SDA output
  io_I2C0SCL_porsccbe,                   // CCBS
  io_I2C0SCL_porsclhsmode,               // SCL high-speed mode select
  io_I2C0SCL_porsclnmode,                // SCL non-I2C mode select
  io_I2C0SCL_porsdhsmode,                // SDA high-speed mode select
  io_I2C0SCL_porsdanmode,                // SDA non-I2C mode select
  io_I2C0SCL_porsdagzn,                  // SDA active-low tri-state and open drain enable

  // I2C1SCL interface
  io_I2C1SCL_piscl,                      // SCL input
  io_I2C1SCL_pisda,                      // SDA input
  io_I2C1SCL_porscl,                     // SCL output
  io_I2C1SCL_porsda,                     // SDA output
  io_I2C1SCL_porsccbe,                   // CCBS
  io_I2C1SCL_porsclhsmode,               // SCL high-speed mode select
  io_I2C1SCL_porsclnmode,                // SCL non-I2C mode select
  io_I2C1SCL_porsdhsmode,                // SDA high-speed mode select
  io_I2C1SCL_porsdanmode,                // SDA non-I2C mode select
  io_I2C1SCL_porsdagzn,                  // SDA active-low tri-state and open drain enable

  // I2C2SCL interface
  io_I2C2SCL_piscl,                      // SCL input
  io_I2C2SCL_pisda,                      // SDA input
  io_I2C2SCL_porscl,                     // SCL output
  io_I2C2SCL_porsda,                     // SDA output
  io_I2C2SCL_porsccbe,                   // CCBS
  io_I2C2SCL_porsclhsmode,               // SCL high-speed mode select
  io_I2C2SCL_porsclnmode,                // SCL non-I2C mode select
  io_I2C2SCL_porsdhsmode,                // SDA high-speed mode select
  io_I2C2SCL_porsdanmode,                // SDA non-I2C mode select
  io_I2C2SCL_porsdagzn,                  // SDA active-low tri-state and open drain enable

  // I2C3SCL interface
  io_I2C3SCL_piscl,                      // SCL input
  io_I2C3SCL_pisda,                      // SDA input
  io_I2C3SCL_porscl,                     // SCL output
  io_I2C3SCL_porsda,                     // SDA output
  io_I2C3SCL_porsccbe,                   // CCBS
  io_I2C3SCL_porsclhsmode,               // SCL high-speed mode select
  io_I2C3SCL_porsclnmode,                // SCL non-I2C mode select
  io_I2C3SCL_porsdhsmode,                // SDA high-speed mode select
  io_I2C3SCL_porsdanmode,                // SDA non-I2C mode select
  io_I2C3SCL_porsdagzn,                  // SDA active-low tri-state and open drain enable

  // XSPI0 interface
  io_XSPI0_mst_in_clk,                   // xspi loopback clock
  io_XSPI0_out_clk,                      // xspi clock out
  io_XSPI0_cs_o,                         // Peripheral Select\n0 - Flash device selected\n1 - Flash device not selected
  io_XSPI0_data_i,                       // Input data from Flash device
  io_XSPI0_data_o,                       // Output Data to flash device
  io_XSPI0_data_oe_n,                    // Flash device output enable\n0 - Enabled\n1 - Not enabled
  io_XSPI0_data_mask_o,                  // Output Data mask needed for Hyperbus protocol
  io_XSPI0_data_mask_oe_n,               // Output Data mask output enable needed for Hyperbus protocol
  io_XSPI0_reset_out,                    // Software controlled separated o/p Hardware Resets for external Flash Devices
  io_XSPI0_reset_in,                     // Software controlled separated i/p Hardware Resets for external Flash Devices
  io_XSPI0_intr_n,                       //  Interrupt input from the Target
  io_XSPI0_dqs_clk,                      // FLASH device DQS

  // CAN0 interface
  io_CAN0_txd,                           // CAN bus Transmit Data
  io_CAN0_rxd,                           // CAN bus Receive Data

  // CAN1 interface
  io_CAN1_txd,                           // CAN bus Transmit Data
  io_CAN1_rxd,                           // CAN bus Receive Data

  // CAN2 interface
  io_CAN2_txd,                           // CAN bus Transmit Data
  io_CAN2_rxd,                           // CAN bus Receive Data

  // CAN3 interface
  io_CAN3_txd,                           // CAN bus Transmit Data
  io_CAN3_rxd,                           // CAN bus Receive Data

  // CAN4 interface
  io_CAN4_txd,                           // CAN bus Transmit Data
  io_CAN4_rxd,                           // CAN bus Receive Data

  // CAN5 interface
  io_CAN5_txd,                           // CAN bus Transmit Data
  io_CAN5_rxd,                           // CAN bus Receive Data

  // CAN6 interface
  io_CAN6_txd,                           // CAN bus Transmit Data
  io_CAN6_rxd,                           // CAN bus Receive Data

  // CAN7 interface
  io_CAN7_txd,                           // CAN bus Transmit Data
  io_CAN7_rxd,                           // CAN bus Receive Data

  // CAN8 interface
  io_CAN8_txd,                           // CAN bus Transmit Data
  io_CAN8_rxd,                           // CAN bus Receive Data

  // CAN9 interface
  io_CAN9_txd,                           // CAN bus Transmit Data
  io_CAN9_rxd,                           // CAN bus Receive Data

  // CAN10 interface
  io_CAN10_txd,                          // CAN bus Transmit Data
  io_CAN10_rxd,                          // CAN bus Receive Data

  // CAN11 interface
  io_CAN11_txd,                          // CAN bus Transmit Data
  io_CAN11_rxd,                          // CAN bus Receive Data

  // LIN0 interface
  io_LIN0_txd,                           // Serial Data Transmission
  io_LIN0_rxd,                           // Serial Data Reception
  io_LIN0_tr_en,                         // Transceiver enable

  // LIN1 interface
  io_LIN1_txd,                           // Serial Data Transmission
  io_LIN1_rxd,                           // Serial Data Reception
  io_LIN1_tr_en,                         // Transceiver enable

  // LIN2 interface
  io_LIN2_txd,                           // Serial Data Transmission
  io_LIN2_rxd,                           // Serial Data Reception
  io_LIN2_tr_en,                         // Transceiver enable

  // LIN3 interface
  io_LIN3_txd,                           // Serial Data Transmission
  io_LIN3_rxd,                           // Serial Data Reception
  io_LIN3_tr_en,                         // Transceiver enable

  // LIN4 interface
  io_LIN4_txd,                           // Serial Data Transmission
  io_LIN4_rxd,                           // Serial Data Reception
  io_LIN4_tr_en,                         // Transceiver enable

  // LIN5 interface
  io_LIN5_txd,                           // Serial Data Transmission
  io_LIN5_rxd,                           // Serial Data Reception
  io_LIN5_tr_en,                         // Transceiver enable

  // LIN6 interface
  io_LIN6_txd,                           // Serial Data Transmission
  io_LIN6_rxd,                           // Serial Data Reception
  io_LIN6_tr_en,                         // Transceiver enable

  // LIN7 interface
  io_LIN7_txd,                           // Serial Data Transmission
  io_LIN7_rxd,                           // Serial Data Reception
  io_LIN7_tr_en,                         // Transceiver enable

  // UART_IO interface
  io_UART0_cd_n,                         
  io_UART0_cts_n,                        
  io_UART0_dsr_n,                        
  io_UART0_dtr_n,                        
  io_UART0_out1,                         
  io_UART0_out2,                         
  io_UART0_ri_n,                         
  io_UART0_rts_n,                        
  io_UART0_rx,                           
  io_UART0_tx,                           

  // UART_IO interface
  io_UART1_cd_n,                         
  io_UART1_cts_n,                        
  io_UART1_dsr_n,                        
  io_UART1_dtr_n,                        
  io_UART1_out1,                         
  io_UART1_out2,                         
  io_UART1_ri_n,                         
  io_UART1_rts_n,                        
  io_UART1_rx,                           
  io_UART1_tx,                           

  // SENT0 interface
  io_SENT0_soc_ext_trig_i,               // SoC external triggers
  io_SENT0_tstamp_val_i,                 // Timestamp value
  io_SENT0_rxd_i,                        // Data input
  io_SENT0_rxd_o,                        // Data output
  io_SENT0_rxd_oen_o,                    // Data output enable

  // SENT1 interface
  io_SENT1_soc_ext_trig_i,               // SoC external triggers
  io_SENT1_tstamp_val_i,                 // Timestamp value
  io_SENT1_rxd_i,                        // Data input
  io_SENT1_rxd_o,                        // Data output
  io_SENT1_rxd_oen_o,                    // Data output enable

  // SENT2 interface
  io_SENT2_soc_ext_trig_i,               // SoC external triggers
  io_SENT2_tstamp_val_i,                 // Timestamp value
  io_SENT2_rxd_i,                        // Data input
  io_SENT2_rxd_o,                        // Data output
  io_SENT2_rxd_oen_o,                    // Data output enable

  // SENT3 interface
  io_SENT3_soc_ext_trig_i,               // SoC external triggers
  io_SENT3_tstamp_val_i,                 // Timestamp value
  io_SENT3_rxd_i,                        // Data input
  io_SENT3_rxd_o,                        // Data output
  io_SENT3_rxd_oen_o,                    // Data output enable

  // SENT4 interface
  io_SENT4_soc_ext_trig_i,               // SoC external triggers
  io_SENT4_tstamp_val_i,                 // Timestamp value
  io_SENT4_rxd_i,                        // Data input
  io_SENT4_rxd_o,                        // Data output
  io_SENT4_rxd_oen_o,                    // Data output enable

  // SENT5 interface
  io_SENT5_soc_ext_trig_i,               // SoC external triggers
  io_SENT5_tstamp_val_i,                 // Timestamp value
  io_SENT5_rxd_i,                        // Data input
  io_SENT5_rxd_o,                        // Data output
  io_SENT5_rxd_oen_o,                    // Data output enable

  // MIBSPI0CLK interface
  io_MIBSPI0CLK_clock,                   // Module/peripheral clock

  // MIBSPI0PICO interface
  io_MIBSPI0PICO_in,                     // Input
  io_MIBSPI0PICO_out,                    // Output
  io_MIBSPI0PICO_oen,                    // Output enable

  // MIBSPI0POCI interface
  io_MIBSPI0POCI_in,                     // Input
  io_MIBSPI0POCI_out,                    // Output
  io_MIBSPI0POCI_oen,                    // Output enable

  // MIBSPI0CS0 interface
  io_MIBSPI0CS0_in,                      // Input
  io_MIBSPI0CS0_out,                     // Output
  io_MIBSPI0CS0_oen,                     // Output enable

  // MIBSPI0CS1 interface
  io_MIBSPI0CS1_in,                      // Input
  io_MIBSPI0CS1_out,                     // Output
  io_MIBSPI0CS1_oen,                     // Output enable

  // MIBSPI0CS2 interface
  io_MIBSPI0CS2_in,                      // Input
  io_MIBSPI0CS2_out,                     // Output
  io_MIBSPI0CS2_oen,                     // Output enable

  // MIBSPI0CS3 interface
  io_MIBSPI0CS3_in,                      // Input
  io_MIBSPI0CS3_out,                     // Output
  io_MIBSPI0CS3_oen,                     // Output enable

  // MIBSPI0CS4 interface
  io_MIBSPI0CS4_in,                      // Input
  io_MIBSPI0CS4_out,                     // Output
  io_MIBSPI0CS4_oen,                     // Output enable

  // MIBSPI0CS5 interface
  io_MIBSPI0CS5_in,                      // Input
  io_MIBSPI0CS5_out,                     // Output
  io_MIBSPI0CS5_oen,                     // Output enable

  // MIBSPI0CS6 interface
  io_MIBSPI0CS6_in,                      // Input
  io_MIBSPI0CS6_out,                     // Output
  io_MIBSPI0CS6_oen,                     // Output enable

  // MIBSPI0CS7 interface
  io_MIBSPI0CS7_in,                      // Input
  io_MIBSPI0CS7_out,                     // Output
  io_MIBSPI0CS7_oen,                     // Output enable

  // MIBSPI0CS8 interface
  io_MIBSPI0CS8_in,                      // Input
  io_MIBSPI0CS8_out,                     // Output
  io_MIBSPI0CS8_oen,                     // Output enable

  // MIBSPI0CS9 interface
  io_MIBSPI0CS9_in,                      // Input
  io_MIBSPI0CS9_out,                     // Output
  io_MIBSPI0CS9_oen,                     // Output enable

  // MIBSPI0CS10 interface
  io_MIBSPI0CS10_in,                     // Input
  io_MIBSPI0CS10_out,                    // Output
  io_MIBSPI0CS10_oen,                    // Output enable

  // MIBSPI0CS11 interface
  io_MIBSPI0CS11_in,                     // Input
  io_MIBSPI0CS11_out,                    // Output
  io_MIBSPI0CS11_oen,                    // Output enable

  // MIBSPI1CLK interface
  io_MIBSPI1CLK_clock,                   // Module/peripheral clock

  // MIBSPI1PICO interface
  io_MIBSPI1PICO_in,                     // Input
  io_MIBSPI1PICO_out,                    // Output
  io_MIBSPI1PICO_oen,                    // Output enable

  // MIBSPI1POCI interface
  io_MIBSPI1POCI_in,                     // Input
  io_MIBSPI1POCI_out,                    // Output
  io_MIBSPI1POCI_oen,                    // Output enable

  // MIBSPI1CS0 interface
  io_MIBSPI1CS0_in,                      // Input
  io_MIBSPI1CS0_out,                     // Output
  io_MIBSPI1CS0_oen,                     // Output enable

  // MIBSPI1CS1 interface
  io_MIBSPI1CS1_in,                      // Input
  io_MIBSPI1CS1_out,                     // Output
  io_MIBSPI1CS1_oen,                     // Output enable

  // MIBSPI1CS2 interface
  io_MIBSPI1CS2_in,                      // Input
  io_MIBSPI1CS2_out,                     // Output
  io_MIBSPI1CS2_oen,                     // Output enable

  // MIBSPI1CS3 interface
  io_MIBSPI1CS3_in,                      // Input
  io_MIBSPI1CS3_out,                     // Output
  io_MIBSPI1CS3_oen,                     // Output enable

  // MIBSPI1CS4 interface
  io_MIBSPI1CS4_in,                      // Input
  io_MIBSPI1CS4_out,                     // Output
  io_MIBSPI1CS4_oen,                     // Output enable

  // MIBSPI1CS5 interface
  io_MIBSPI1CS5_in,                      // Input
  io_MIBSPI1CS5_out,                     // Output
  io_MIBSPI1CS5_oen,                     // Output enable

  // MIBSPI1CS6 interface
  io_MIBSPI1CS6_in,                      // Input
  io_MIBSPI1CS6_out,                     // Output
  io_MIBSPI1CS6_oen,                     // Output enable

  // MIBSPI1CS7 interface
  io_MIBSPI1CS7_in,                      // Input
  io_MIBSPI1CS7_out,                     // Output
  io_MIBSPI1CS7_oen,                     // Output enable

  // MIBSPI1CS8 interface
  io_MIBSPI1CS8_in,                      // Input
  io_MIBSPI1CS8_out,                     // Output
  io_MIBSPI1CS8_oen,                     // Output enable

  // MIBSPI1CS9 interface
  io_MIBSPI1CS9_in,                      // Input
  io_MIBSPI1CS9_out,                     // Output
  io_MIBSPI1CS9_oen,                     // Output enable

  // MIBSPI1CS10 interface
  io_MIBSPI1CS10_in,                     // Input
  io_MIBSPI1CS10_out,                    // Output
  io_MIBSPI1CS10_oen,                    // Output enable

  // MIBSPI1CS11 interface
  io_MIBSPI1CS11_in,                     // Input
  io_MIBSPI1CS11_out,                    // Output
  io_MIBSPI1CS11_oen,                    // Output enable

  // SPI2CLK interface
  io_SPI2CLK_clock,                      // Module/peripheral clock

  // SPI2PICO interface
  io_SPI2PICO_in,                        // Input
  io_SPI2PICO_out,                       // Output
  io_SPI2PICO_oen,                       // Output enable

  // SPI2POCI interface
  io_SPI2POCI_in,                        // Input
  io_SPI2POCI_out,                       // Output
  io_SPI2POCI_oen,                       // Output enable

  // SPI2CS0 interface
  io_SPI2CS0_in,                         // Input
  io_SPI2CS0_out,                        // Output
  io_SPI2CS0_oen,                        // Output enable

  // SPI2CS1 interface
  io_SPI2CS1_in,                         // Input
  io_SPI2CS1_out,                        // Output
  io_SPI2CS1_oen,                        // Output enable

  // SPI2CS2 interface
  io_SPI2CS2_in,                         // Input
  io_SPI2CS2_out,                        // Output
  io_SPI2CS2_oen,                        // Output enable

  // SPI2CS3 interface
  io_SPI2CS3_in,                         // Input
  io_SPI2CS3_out,                        // Output
  io_SPI2CS3_oen,                        // Output enable

  // SPI2CS4 interface
  io_SPI2CS4_in,                         // Input
  io_SPI2CS4_out,                        // Output
  io_SPI2CS4_oen,                        // Output enable

  // SPI2CS5 interface
  io_SPI2CS5_in,                         // Input
  io_SPI2CS5_out,                        // Output
  io_SPI2CS5_oen,                        // Output enable

  // SPI3CLK interface
  io_SPI3CLK_clock,                      // Module/peripheral clock

  // SPI3PICO interface
  io_SPI3PICO_in,                        // Input
  io_SPI3PICO_out,                       // Output
  io_SPI3PICO_oen,                       // Output enable

  // SPI3POCI interface
  io_SPI3POCI_in,                        // Input
  io_SPI3POCI_out,                       // Output
  io_SPI3POCI_oen,                       // Output enable

  // SPI3CS0 interface
  io_SPI3CS0_in,                         // Input
  io_SPI3CS0_out,                        // Output
  io_SPI3CS0_oen,                        // Output enable

  // SPI3CS1 interface
  io_SPI3CS1_in,                         // Input
  io_SPI3CS1_out,                        // Output
  io_SPI3CS1_oen,                        // Output enable

  // SPI3CS2 interface
  io_SPI3CS2_in,                         // Input
  io_SPI3CS2_out,                        // Output
  io_SPI3CS2_oen,                        // Output enable

  // SPI3CS3 interface
  io_SPI3CS3_in,                         // Input
  io_SPI3CS3_out,                        // Output
  io_SPI3CS3_oen,                        // Output enable

  // SPI3CS4 interface
  io_SPI3CS4_in,                         // Input
  io_SPI3CS4_out,                        // Output
  io_SPI3CS4_oen,                        // Output enable

  // SPI3CS5 interface
  io_SPI3CS5_in,                         // Input
  io_SPI3CS5_out,                        // Output
  io_SPI3CS5_oen,                        // Output enable

  // SPI4CLK interface
  io_SPI4CLK_clock,                      // Module/peripheral clock

  // SPI4PICO interface
  io_SPI4PICO_in,                        // Input
  io_SPI4PICO_out,                       // Output
  io_SPI4PICO_oen,                       // Output enable

  // SPI4POCI interface
  io_SPI4POCI_in,                        // Input
  io_SPI4POCI_out,                       // Output
  io_SPI4POCI_oen,                       // Output enable

  // SPI4CS0 interface
  io_SPI4CS0_in,                         // Input
  io_SPI4CS0_out,                        // Output
  io_SPI4CS0_oen,                        // Output enable

  // SPI4CS1 interface
  io_SPI4CS1_in,                         // Input
  io_SPI4CS1_out,                        // Output
  io_SPI4CS1_oen,                        // Output enable

  // SPI4CS2 interface
  io_SPI4CS2_in,                         // Input
  io_SPI4CS2_out,                        // Output
  io_SPI4CS2_oen,                        // Output enable

  // SPI4CS3 interface
  io_SPI4CS3_in,                         // Input
  io_SPI4CS3_out,                        // Output
  io_SPI4CS3_oen,                        // Output enable

  // SPI4CS4 interface
  io_SPI4CS4_in,                         // Input
  io_SPI4CS4_out,                        // Output
  io_SPI4CS4_oen,                        // Output enable

  // SPI4CS5 interface
  io_SPI4CS5_in,                         // Input
  io_SPI4CS5_out,                        // Output
  io_SPI4CS5_oen,                        // Output enable

  // SPI5CLK interface
  io_SPI5CLK_clock,                      // Module/peripheral clock

  // SPI5PICO interface
  io_SPI5PICO_in,                        // Input
  io_SPI5PICO_out,                       // Output
  io_SPI5PICO_oen,                       // Output enable

  // SPI5POCI interface
  io_SPI5POCI_in,                        // Input
  io_SPI5POCI_out,                       // Output
  io_SPI5POCI_oen,                       // Output enable

  // SPI5CS0 interface
  io_SPI5CS0_in,                         // Input
  io_SPI5CS0_out,                        // Output
  io_SPI5CS0_oen,                        // Output enable

  // SPI5CS1 interface
  io_SPI5CS1_in,                         // Input
  io_SPI5CS1_out,                        // Output
  io_SPI5CS1_oen,                        // Output enable

  // SPI5CS2 interface
  io_SPI5CS2_in,                         // Input
  io_SPI5CS2_out,                        // Output
  io_SPI5CS2_oen,                        // Output enable

  // SPI5CS3 interface
  io_SPI5CS3_in,                         // Input
  io_SPI5CS3_out,                        // Output
  io_SPI5CS3_oen,                        // Output enable

  // SPI5CS4 interface
  io_SPI5CS4_in,                         // Input
  io_SPI5CS4_out,                        // Output
  io_SPI5CS4_oen,                        // Output enable

  // SPI5CS5 interface
  io_SPI5CS5_in,                         // Input
  io_SPI5CS5_out,                        // Output
  io_SPI5CS5_oen,                        // Output enable

  // SPI6CLK interface
  io_SPI6CLK_clock,                      // Module/peripheral clock

  // SPI6PICO interface
  io_SPI6PICO_in,                        // Input
  io_SPI6PICO_out,                       // Output
  io_SPI6PICO_oen,                       // Output enable

  // SPI6POCI interface
  io_SPI6POCI_in,                        // Input
  io_SPI6POCI_out,                       // Output
  io_SPI6POCI_oen,                       // Output enable

  // SPI6CS0 interface
  io_SPI6CS0_in,                         // Input
  io_SPI6CS0_out,                        // Output
  io_SPI6CS0_oen,                        // Output enable

  // SPI6CS1 interface
  io_SPI6CS1_in,                         // Input
  io_SPI6CS1_out,                        // Output
  io_SPI6CS1_oen,                        // Output enable

  // SPI6CS2 interface
  io_SPI6CS2_in,                         // Input
  io_SPI6CS2_out,                        // Output
  io_SPI6CS2_oen,                        // Output enable

  // SPI6CS3 interface
  io_SPI6CS3_in,                         // Input
  io_SPI6CS3_out,                        // Output
  io_SPI6CS3_oen,                        // Output enable

  // SPI6CS4 interface
  io_SPI6CS4_in,                         // Input
  io_SPI6CS4_out,                        // Output
  io_SPI6CS4_oen,                        // Output enable

  // SPI6CS5 interface
  io_SPI6CS5_in,                         // Input
  io_SPI6CS5_out,                        // Output
  io_SPI6CS5_oen,                        // Output enable

  // SPI7CLK interface
  io_SPI7CLK_clock,                      // Module/peripheral clock

  // SPI7PICO interface
  io_SPI7PICO_in,                        // Input
  io_SPI7PICO_out,                       // Output
  io_SPI7PICO_oen,                       // Output enable

  // SPI7POCI interface
  io_SPI7POCI_in,                        // Input
  io_SPI7POCI_out,                       // Output
  io_SPI7POCI_oen,                       // Output enable

  // SPI7CS0 interface
  io_SPI7CS0_in,                         // Input
  io_SPI7CS0_out,                        // Output
  io_SPI7CS0_oen,                        // Output enable

  // SPI7CS1 interface
  io_SPI7CS1_in,                         // Input
  io_SPI7CS1_out,                        // Output
  io_SPI7CS1_oen,                        // Output enable

  // SPI7CS2 interface
  io_SPI7CS2_in,                         // Input
  io_SPI7CS2_out,                        // Output
  io_SPI7CS2_oen,                        // Output enable

  // SPI7CS3 interface
  io_SPI7CS3_in,                         // Input
  io_SPI7CS3_out,                        // Output
  io_SPI7CS3_oen,                        // Output enable

  // SPI7CS4 interface
  io_SPI7CS4_in,                         // Input
  io_SPI7CS4_out,                        // Output
  io_SPI7CS4_oen,                        // Output enable

  // SPI7CS5 interface
  io_SPI7CS5_in,                         // Input
  io_SPI7CS5_out,                        // Output
  io_SPI7CS5_oen,                        // Output enable

  // SPI8CLK interface
  io_SPI8CLK_clock,                      // Module/peripheral clock

  // SPI8PICO interface
  io_SPI8PICO_in,                        // Input
  io_SPI8PICO_out,                       // Output
  io_SPI8PICO_oen,                       // Output enable

  // SPI8POCI interface
  io_SPI8POCI_in,                        // Input
  io_SPI8POCI_out,                       // Output
  io_SPI8POCI_oen,                       // Output enable

  // SPI8CS0 interface
  io_SPI8CS0_in,                         // Input
  io_SPI8CS0_out,                        // Output
  io_SPI8CS0_oen,                        // Output enable

  // SPI8CS1 interface
  io_SPI8CS1_in,                         // Input
  io_SPI8CS1_out,                        // Output
  io_SPI8CS1_oen,                        // Output enable

  // SPI8CS2 interface
  io_SPI8CS2_in,                         // Input
  io_SPI8CS2_out,                        // Output
  io_SPI8CS2_oen,                        // Output enable

  // SPI8CS3 interface
  io_SPI8CS3_in,                         // Input
  io_SPI8CS3_out,                        // Output
  io_SPI8CS3_oen,                        // Output enable

  // SPI8CS4 interface
  io_SPI8CS4_in,                         // Input
  io_SPI8CS4_out,                        // Output
  io_SPI8CS4_oen,                        // Output enable

  // SPI8CS5 interface
  io_SPI8CS5_in,                         // Input
  io_SPI8CS5_out,                        // Output
  io_SPI8CS5_oen,                        // Output enable

  // SPI9CLK interface
  io_SPI9CLK_clock,                      // Module/peripheral clock

  // SPI9PICO interface
  io_SPI9PICO_in,                        // Input
  io_SPI9PICO_out,                       // Output
  io_SPI9PICO_oen,                       // Output enable

  // SPI9POCI interface
  io_SPI9POCI_in,                        // Input
  io_SPI9POCI_out,                       // Output
  io_SPI9POCI_oen,                       // Output enable

  // SPI9CS0 interface
  io_SPI9CS0_in,                         // Input
  io_SPI9CS0_out,                        // Output
  io_SPI9CS0_oen,                        // Output enable

  // SPI9CS1 interface
  io_SPI9CS1_in,                         // Input
  io_SPI9CS1_out,                        // Output
  io_SPI9CS1_oen,                        // Output enable

  // SPI9CS2 interface
  io_SPI9CS2_in,                         // Input
  io_SPI9CS2_out,                        // Output
  io_SPI9CS2_oen,                        // Output enable

  // SPI9CS3 interface
  io_SPI9CS3_in,                         // Input
  io_SPI9CS3_out,                        // Output
  io_SPI9CS3_oen,                        // Output enable

  // SPI9CS4 interface
  io_SPI9CS4_in,                         // Input
  io_SPI9CS4_out,                        // Output
  io_SPI9CS4_oen,                        // Output enable

  // SPI9CS5 interface
  io_SPI9CS5_in,                         // Input
  io_SPI9CS5_out,                        // Output
  io_SPI9CS5_oen,                        // Output enable

  // PSI5_IO interface
  io_PSI5_0_tx,                          // Serial Data Transmission
  io_PSI5_0_rx,                          // Serial Data Reception

  // PSI5_IO interface
  io_PSI5_1_tx,                          // Serial Data Transmission
  io_PSI5_1_rx,                          // Serial Data Reception

  // PSI5_IO interface
  io_PSI5_2_tx,                          // Serial Data Transmission
  io_PSI5_2_rx,                          // Serial Data Reception

  // PSI5_IO interface
  io_PSI5_3_tx,                          // Serial Data Transmission
  io_PSI5_3_rx                           // Serial Data Reception
);

// Default Interface

// IO PORT
inout             AP0_IO;

// IO PORT
inout             AP1_IO;

// IO PORT
inout             AP10_IO;

// IO PORT
inout             AP11_IO;

// IO PORT
inout             AP12_IO;

// IO PORT
inout             AP13_IO;

// IO PORT
inout             AP14_IO;

// IO PORT
inout             AP15_IO;

// IO PORT
inout             AP16_IO;

// IO PORT
inout             AP17_IO;

// IO PORT
inout             AP18_IO;

// IO PORT
inout             AP19_IO;

// IO PORT
inout             AP2_IO;

// IO PORT
inout             AP20_IO;

// IO PORT
inout             AP21_IO;

// IO PORT
inout             AP22_IO;

// IO PORT
inout             AP23_IO;

// IO PORT
inout             AP24_IO;

// IO PORT
inout             AP25_IO;

// IO PORT
inout             AP26_IO;

// IO PORT
inout             AP27_IO;

// IO PORT
inout             AP28_IO;

// IO PORT
inout             AP29_IO;

// IO PORT
inout             AP3_IO;

// IO PORT
inout             AP30_IO;

// IO PORT
inout             AP31_IO;

// IO PORT
inout             AP32_IO;

// IO PORT
inout             AP33_IO;

// IO PORT
inout             AP34_IO;

// IO PORT
inout             AP35_IO;

// IO PORT
inout             AP36_IO;

// IO PORT
inout             AP37_IO;

// IO PORT
inout             AP38_IO;

// IO PORT
inout             AP39_IO;

// IO PORT
inout             AP4_IO;

// IO PORT
inout             AP40_IO;

// IO PORT
inout             AP41_IO;

// IO PORT
inout             AP42_IO;

// IO PORT
inout             AP43_IO;

// IO PORT
inout             AP44_IO;

// IO PORT
inout             AP45_IO;

// IO PORT
inout             AP46_IO;

// IO PORT
inout             AP47_IO;

// IO PORT
inout             AP5_IO;

// IO PORT
inout             AP6_IO;

// IO PORT
inout             AP7_IO;

// IO PORT
inout             AP8_IO;

// IO PORT
inout             AP9_IO;

// IO PORT
inout             AURORACLKN_IO;

// IO PORT
inout             AURORACLKP_IO;

// IO PORT
inout             AURORADN_IO;

// IO PORT
inout             AURORADP_IO;

// IO PORT
inout             DCDCNMOS_IO;

// IO PORT
inout             DCDCPMOS_IO;

// IO PORT
inout             DP0_0_IO;

// IO PORT
inout             DP0_1_IO;

// IO PORT
inout             DP0_2_IO;

// IO PORT
inout             DP0_3_IO;

// IO PORT
inout             DP0_4_IO;

// IO PORT
inout             DP0_5_IO;

// IO PORT
inout             DP0_6_IO;

// IO PORT
inout             DP0_7_IO;

// IO PORT
inout             DP0_8_IO;

// IO PORT
inout             DP0_9_IO;

// IO PORT
inout             DP0_10_IO;

// IO PORT
inout             DP0_11_IO;

// IO PORT
inout             DP0_12_IO;

// IO PORT
inout             DP0_13_IO;

// IO PORT
inout             DP0_14_IO;

// IO PORT
inout             DP0_15_IO;

// IO PORT
inout             DP0_16_IO;

// IO PORT
inout             DP0_17_IO;

// IO PORT
inout             DP0_18_IO;

// IO PORT
inout             DP0_19_IO;

// IO PORT
inout             DP0_20_IO;

// IO PORT
inout             DP0_21_IO;

// IO PORT
inout             DP0_22_IO;

// IO PORT
inout             DP0_23_IO;

// IO PORT
inout             DP0_24_IO;

// IO PORT
inout             DP0_25_IO;

// IO PORT
inout             DP0_26_IO;

// IO PORT
inout             DP0_27_IO;

// IO PORT
inout             DP0_28_IO;

// IO PORT
inout             DP0_29_IO;

// IO PORT
inout             DP0_30_IO;

// IO PORT
inout             DP0_31_IO;

// IO PORT
inout             DP1_0_IO;

// IO PORT
inout             DP1_1_IO;

// IO PORT
inout             DP1_2_IO;

// IO PORT
inout             DP1_3_IO;

// IO PORT
inout             DP1_4_IO;

// IO PORT
inout             DP1_5_IO;

// IO PORT
inout             DP1_6_IO;

// IO PORT
inout             DP1_7_IO;

// IO PORT
inout             DP1_8_IO;

// IO PORT
inout             DP1_9_IO;

// IO PORT
inout             DP1_10_IO;

// IO PORT
inout             DP1_11_IO;

// IO PORT
inout             DP1_12_IO;

// IO PORT
inout             DP1_13_IO;

// IO PORT
inout             DP1_14_IO;

// IO PORT
inout             DP1_15_IO;

// IO PORT
inout             DP1_16_IO;

// IO PORT
inout             DP1_17_IO;

// IO PORT
inout             DP1_18_IO;

// IO PORT
inout             DP1_19_IO;

// IO PORT
inout             DP1_20_IO;

// IO PORT
inout             DP1_21_IO;

// IO PORT
inout             DP1_22_IO;

// IO PORT
inout             DP1_23_IO;

// IO PORT
inout             DP1_24_IO;

// IO PORT
inout             DP1_25_IO;

// IO PORT
inout             DP1_26_IO;

// IO PORT
inout             DP1_27_IO;

// IO PORT
inout             DP1_28_IO;

// IO PORT
inout             DP1_29_IO;

// IO PORT
inout             DP1_30_IO;

// IO PORT
inout             DP1_31_IO;

// IO PORT
inout             DP2_0_IO;

// IO PORT
inout             DP2_1_IO;

// IO PORT
inout             DP2_2_IO;

// IO PORT
inout             DP2_3_IO;

// IO PORT
inout             DP2_4_IO;

// IO PORT
inout             DP2_5_IO;

// IO PORT
inout             DP2_6_IO;

// IO PORT
inout             DP2_7_IO;

// IO PORT
inout             DP2_8_IO;

// IO PORT
inout             DP2_9_IO;

// IO PORT
inout             DP2_10_IO;

// IO PORT
inout             DP2_11_IO;

// IO PORT
inout             DP2_12_IO;

// IO PORT
inout             DP2_13_IO;

// IO PORT
inout             DP2_14_IO;

// IO PORT
inout             DP2_15_IO;

// IO PORT
inout             DP2_16_IO;

// IO PORT
inout             DP2_17_IO;

// IO PORT
inout             DP2_18_IO;

// IO PORT
inout             DP2_19_IO;

// IO PORT
inout             DP2_20_IO;

// IO PORT
inout             DP2_21_IO;

// IO PORT
inout             DP2_22_IO;

// IO PORT
inout             DP2_23_IO;

// IO PORT
inout             DP2_24_IO;

// IO PORT
inout             DP2_25_IO;

// IO PORT
inout             DP2_26_IO;

// IO PORT
inout             DP2_27_IO;

// IO PORT
inout             DP2_28_IO;

// IO PORT
inout             DP2_29_IO;

// IO PORT
inout             DP2_30_IO;

// IO PORT
inout             DP2_31_IO;

// IO PORT
inout             DP3_0_IO;

// IO PORT
inout             DP3_1_IO;

// IO PORT
inout             DP3_2_IO;

// IO PORT
inout             DP3_3_IO;

// IO PORT
inout             DP3_4_IO;

// IO PORT
inout             DP3_5_IO;

// IO PORT
inout             DP3_6_IO;

// IO PORT
inout             DP3_7_IO;

// IO PORT
inout             DP3_8_IO;

// IO PORT
inout             DP3_9_IO;

// IO PORT
inout             DP3_10_IO;

// IO PORT
inout             DP3_11_IO;

// IO PORT
inout             DP3_12_IO;

// IO PORT
inout             DP3_13_IO;

// IO PORT
inout             DP3_14_IO;

// IO PORT
inout             DP3_15_IO;

// IO PORT
inout             DP3_16_IO;

// IO PORT
inout             DP3_17_IO;

// IO PORT
inout             DP3_18_IO;

// IO PORT
inout             DP3_19_IO;

// IO PORT
inout             DP3_20_IO;

// IO PORT
inout             DP3_21_IO;

// IO PORT
inout             DP3_22_IO;

// IO PORT
inout             DP3_23_IO;

// IO PORT
inout             DP3_24_IO;

// IO PORT
inout             DP3_25_IO;

// IO PORT
inout             DP3_26_IO;

// IO PORT
inout             DP3_27_IO;

// IO PORT
inout             DP3_28_IO;

// IO PORT
inout             DP3_29_IO;

// IO PORT
inout             DP3_30_IO;

// IO PORT
inout             DP3_31_IO;

// IO PORT
inout             DP4_0_IO;

// IO PORT
inout             DP4_1_IO;

// IO PORT
inout             DP4_2_IO;

// IO PORT
inout             DP4_3_IO;

// IO PORT
inout             DP4_4_IO;

// IO PORT
inout             DP4_5_IO;

// IO PORT
inout             DP4_6_IO;

// IO PORT
inout             DP4_7_IO;

// IO PORT
inout             DP4_8_IO;

// IO PORT
inout             DP4_9_IO;

// IO PORT
inout             DP4_10_IO;

// IO PORT
inout             DP4_11_IO;

// IO PORT
inout             DP4_12_IO;

// IO PORT
inout             DP4_13_IO;

// IO PORT
inout             DP4_14_IO;

// IO PORT
inout             DP4_15_IO;

// IO PORT
inout             DP4_16_IO;

// IO PORT
inout             DP4_17_IO;

// IO PORT
inout             DP4_18_IO;

// IO PORT
inout             DP4_19_IO;

// IO PORT
inout             DP4_20_IO;

// IO PORT
inout             DP4_21_IO;

// IO PORT
inout             DP4_22_IO;

// IO PORT
inout             DP4_23_IO;

// IO PORT
inout             DP4_24_IO;

// IO PORT
inout             DP4_25_IO;

// IO PORT
inout             DP4_26_IO;

// IO PORT
inout             DP4_27_IO;

// IO PORT
inout             DP4_28_IO;

// IO PORT
inout             DP4_29_IO;

// IO PORT
inout             DP4_30_IO;

// IO PORT
inout             DP4_31_IO;

// IO PORT
inout             DP5_0_IO;

// IO PORT
inout             DP5_1_IO;

// IO PORT
inout             DP5_2_IO;

// IO PORT
inout             DP5_3_IO;

// IO PORT
inout             DP5_4_IO;

// IO PORT
inout             DP5_5_IO;

// IO PORT
inout             DP5_6_IO;

// IO PORT
inout             DP5_7_IO;

// IO PORT
inout             DP5_8_IO;

// IO PORT
inout             DP5_9_IO;

// IO PORT
inout             DP5_10_IO;

// IO PORT
inout             DP5_11_IO;

// IO PORT
inout             DP5_12_IO;

// IO PORT
inout             DP5_13_IO;

// IO PORT
inout             DP5_14_IO;

// IO PORT
inout             DP5_15_IO;

// IO PORT
inout             DP5_16_IO;

// IO PORT
inout             DP5_17_IO;

// IO PORT
inout             DP5_18_IO;

// IO PORT
inout             DP5_19_IO;

// IO PORT
inout             DP5_20_IO;

// IO PORT
inout             DP5_21_IO;

// IO PORT
inout             DP5_22_IO;

// IO PORT
inout             DP5_23_IO;

// IO PORT
inout             DP5_24_IO;

// IO PORT
inout             DP5_25_IO;

// IO PORT
inout             DP5_26_IO;

// IO PORT
inout             DP5_27_IO;

// IO PORT
inout             DP5_28_IO;

// IO PORT
inout             DP5_29_IO;

// IO PORT
inout             DP5_30_IO;

// IO PORT
inout             DP5_31_IO;

// IO PORT
inout             DP6_0_IO;

// IO PORT
inout             DP6_1_IO;

// IO PORT
inout             DP6_2_IO;

// IO PORT
inout             DP6_3_IO;

// IO PORT
inout             DP6_4_IO;

// IO PORT
inout             DP6_5_IO;

// IO PORT
inout             DP6_6_IO;

// IO PORT
inout             DP6_7_IO;

// IO PORT
inout             DP6_8_IO;

// IO PORT
inout             DP6_9_IO;

// IO PORT
inout             DP6_10_IO;

// IO PORT
inout             DP6_11_IO;

// IO PORT
inout             DP6_12_IO;

// IO PORT
inout             DP6_13_IO;

// IO PORT
inout             DP6_14_IO;

// IO PORT
inout             DP6_15_IO;

// IO PORT
inout             DP6_16_IO;

// IO PORT
inout             DP6_17_IO;

// IO PORT
inout             DP6_18_IO;

// IO PORT
inout             DP6_19_IO;

// IO PORT
inout             DP6_20_IO;

// IO PORT
inout             DP6_21_IO;

// IO PORT
inout             DP6_22_IO;

// IO PORT
inout             DP6_23_IO;

// IO PORT
inout             DP6_24_IO;

// IO PORT
inout             DP6_25_IO;

// IO PORT
inout             DP6_26_IO;

// IO PORT
inout             DP6_27_IO;

// IO PORT
inout             DP7_0_IO;

// IO PORT
inout             DP7_1_IO;

// IO PORT
inout             DP7_2_IO;

// IO PORT
inout             DP7_3_IO;

// IO PORT
inout             DP7_4_IO;

// IO PORT
inout             DP7_5_IO;

// IO PORT
inout             DP7_6_IO;

// IO PORT
inout             DP7_7_IO;

// IO PORT
inout             DP7_8_IO;

// IO PORT
inout             DP7_9_IO;

// IO PORT
inout             DP7_10_IO;

// IO PORT
inout             DP7_11_IO;

// IO PORT
inout             DP7_12_IO;

// IO PORT
inout             DP7_13_IO;

// IO PORT
inout             DP7_14_IO;

// IO PORT
inout             DP7_15_IO;

// IO PORT
inout             ERROR_IO;

// IO PORT
inout             EXTPMICEN_IO;

// IO PORT
inout             FLASHTESTPAD1FT_IO;

// IO PORT
inout             FLASHTESTPAD2_IO;

// IO PORT
inout             FLASHTESTPAD3FT_IO;

// IO PORT
inout             FLASHTESTPAD4_IO;

// IO PORT
inout             FLASHTESTPAD5_IO;

// IO PORT
inout             MP0_0_IO;

// IO PORT
inout             MP0_1_IO;

// IO PORT
inout             MP0_2_IO;

// IO PORT
inout             MP0_3_IO;

// IO PORT
inout             MP0_4_IO;

// IO PORT
inout             MP0_5_IO;

// IO PORT
inout             MP0_6_IO;

// IO PORT
inout             MP0_7_IO;

// IO PORT
inout             MP0_8_IO;

// IO PORT
inout             MP0_9_IO;

// IO PORT
inout             MP0_10_IO;

// IO PORT
inout             MP0_11_IO;

// IO PORT
inout             MP0_12_IO;

// IO PORT
inout             MP0_13_IO;

// IO PORT
inout             MP0_14_IO;

// IO PORT
inout             MP0_15_IO;

// IO PORT
inout             MP0_16_IO;

// IO PORT
inout             MP0_17_IO;

// IO PORT
inout             MP0_18_IO;

// IO PORT
inout             MP0_19_IO;

// IO PORT
inout             MP0_20_IO;

// IO PORT
inout             MP0_21_IO;

// IO PORT
inout             MP0_22_IO;

// IO PORT
inout             MP0_23_IO;

// IO PORT
inout             MP0_24_IO;

// IO PORT
inout             MP0_25_IO;

// IO PORT
inout             MP0_26_IO;

// IO PORT
inout             MP0_27_IO;

// IO PORT
inout             MP0_28_IO;

// IO PORT
inout             MP0_29_IO;

// IO PORT
inout             MP0_30_IO;

// IO PORT
inout             MP0_31_IO;

// IO PORT
inout             MP1_0_IO;

// IO PORT
inout             MP1_1_IO;

// IO PORT
inout             MP1_2_IO;

// IO PORT
inout             MP1_3_IO;

// IO PORT
inout             MP1_4_IO;

// IO PORT
inout             MP1_5_IO;

// IO PORT
inout             MP1_6_IO;

// IO PORT
inout             MP1_7_IO;

// IO PORT
inout             MP1_8_IO;

// IO PORT
inout             MP1_9_IO;

// IO PORT
inout             MP1_10_IO;

// IO PORT
inout             MP1_11_IO;

// IO PORT
inout             MP1_12_IO;

// IO PORT
inout             MP1_13_IO;

// IO PORT
inout             MP1_14_IO;

// IO PORT
inout             MP1_15_IO;

// IO PORT
inout             MP2_0_IO;

// IO PORT
inout             MP2_1_IO;

// IO PORT
inout             MP2_2_IO;

// IO PORT
inout             MP2_3_IO;

// IO PORT
inout             MP2_4_IO;

// IO PORT
inout             MP2_5_IO;

// IO PORT
inout             MP2_6_IO;

// IO PORT
inout             MP2_7_IO;

// IO PORT
inout             MP2_8_IO;

// IO PORT
inout             MP2_9_IO;

// IO PORT
inout             MP2_10_IO;

// IO PORT
inout             MP2_11_IO;

// IO PORT
inout             MP2_12_IO;

// IO PORT
inout             MP2_13_IO;

// IO PORT
inout             MP2_14_IO;

// IO PORT
inout             MP2_15_IO;

// IO PORT
inout             PWR_ON_RSTn_IO;

// IO PORT
inout             RESETOUTn_IO;

// IO PORT
inout             SGMII0RXN_IO;

// IO PORT
inout             SGMII0RXP_IO;

// IO PORT
inout             SGMII0TXN_IO;

// IO PORT
inout             SGMII0TXP_IO;

// IO PORT
inout             SGMII1RXN_IO;

// IO PORT
inout             SGMII1RXP_IO;

// IO PORT
inout             SGMII1TXN_IO;

// IO PORT
inout             SGMII1TXP_IO;

// IO PORT
inout             SGMII2RXN_IO;

// IO PORT
inout             SGMII2RXP_IO;

// IO PORT
inout             SGMII2TXN_IO;

// IO PORT
inout             SGMII2TXP_IO;

// IO PORT
inout             SPI0LPBCLKUNB_IO;

// IO PORT
inout             SPI1LPBCLKUNB_IO;

// IO PORT
inout             SPI2LPBCLKUNB_IO;

// IO PORT
inout             SPI3LPBCLKUNB_IO;

// IO PORT
inout             SPI4LPBCLKUNB_IO;

// IO PORT
inout             SPI5LPBCLKUNB_IO;

// IO PORT
inout             SPI6LPBCLKUNB_IO;

// IO PORT
inout             SPI7LPBCLKUNB_IO;

// IO PORT
inout             SPI8LPBCLKUNB_IO;

// IO PORT
inout             SPI9LPBCLKUNB_IO;

// IO PORT
inout             TCK_IO;

// IO PORT
inout             TDI_IO;

// IO PORT
inout             TDO_IO;

// IO PORT
inout             TMS_IO;

// IO PORT
inout             TRSTN_IO;

// IO PORT
inout             VDDS_REF_LPD_HI_IO;

// IO PORT
inout             VDDS_REF_LPD_LO_IO;

// IO PORT
inout             VDDS_REF_SD_HI_IO;

// IO PORT
inout             VDDS_REF_SD_LO_IO;

// IO PORT
inout             VDDS_REF0_HI_IO;

// IO PORT
inout             VDDS_REF0_LO_IO;

// IO PORT
inout             VDDS_REF1_HI_IO;

// IO PORT
inout             VDDS_REF1_LO_IO;

// IO PORT
inout             VDDS_REF2_HI_IO;

// IO PORT
inout             VDDS_REF2_LO_IO;

// IO PORT
inout             X1_IO;

// IO PORT
inout             X2_IO;

// IO PORT
inout             XSPI0LBCLKUNB_IO;

// PINMUX Clock interface
input             pinmux_clock;

// PINMUX Reset interface
input             pinmux_reset_n;

// GPIO Clock interface
input             gpio_clock;

// IO Clock interface
input             io_clock;

// IO Reset interface
input             gpio_reset_n;

// System Reset interface
input             sys_reset_n;

// IO Reset interface
input             io_reset_n;

// Clock Interface
input             xbar_clk_clock;

// Reset Interface
input             xbar_rst_reset_n;

// jtag_interface
output            jtag_tck;
output            jtag_trst_n;
output            jtag_tdi;
output            jtag_tms;
input             jtag_tdo_oe_n;
input             jtag_tdo;

// o_xrsn_pm_b_reset  interface
output            o_xrsn_pm_b_reset_n;

// o_xrsn_sw_fast_reset  interface
output            o_xrsn_sw_fast_reset_n;

// o_porsn_frompmm_pm_d_reset  interface
output            o_porsn_frompmm_pm_d_reset_n;

// o_porsn_pm_b_reset  interface
output            o_porsn_pm_b_reset_n;

// o_porsn_sw_pm_a_reset  interface
output            o_porsn_sw_pm_a_reset_n;

// o_porsn_sw_pm_b_reset  interface
output            o_porsn_sw_pm_b_reset_n;

// o_porsn_sw_pm_d_reset  interface
output            o_porsn_sw_pm_d_reset_n;

// o_porsn_frompad_reset  interface
output            o_porsn_frompad_reset_n;

// o_porsn_frompmm_pm_a_reset  interface
output            o_porsn_frompmm_pm_a_reset_n;

// o_porsn_sw_streched_pm_a_reset  interface
output            o_porsn_sw_streched_pm_a_reset_n;

// o_porsn_frompmm_pm_b_reset  interface
output            o_porsn_frompmm_pm_b_reset_n;

// o_porsn_sw_streched_pm_b_reset  interface
output            o_porsn_sw_streched_pm_b_reset_n;

// o_xrsn_frompad_reset  interface
output            o_xrsn_frompad_reset_n;

// o_xrsn_sw_streched_reset  interface
output            o_xrsn_sw_streched_reset_n;

// CBA_VBUSP_4_0 BUS Slave view interface
input       [11:0] io_vbusp_slv_routeid;
input       [11:0] io_vbusp_slv_xid;
input             io_vbusp_slv_req;
input             io_vbusp_slv_dir;
input       [31:0] io_vbusp_slv_address;
input        [2:0] io_vbusp_slv_xcnt;
input        [3:0] io_vbusp_slv_byten;
input       [31:0] io_vbusp_slv_wdata;
output            io_vbusp_slv_wready;
output      [31:0] io_vbusp_slv_rdatap;
output       [2:0] io_vbusp_slv_rstatus;
output            io_vbusp_slv_rready;
input        [1:0] io_vbusp_slv_dtype;
input        [1:0] io_vbusp_slv_priv;
input        [7:0] io_vbusp_slv_privid;
input             io_vbusp_slv_secure;
input             io_vbusp_slv_emudbg;

// LPD_CAN0TX interface
input             io_LPD_CAN0TX_txd;
output            io_LPD_CAN0TX_rxd;

// LPD_CAN0RX interface
input             io_LPD_CAN0RX_txd;
output            io_LPD_CAN0RX_rxd;

// LPD_LIN0TX interface
input             io_LPD_LIN0TX_txd;
output            io_LPD_LIN0TX_rxd;
input             io_LPD_LIN0TX_tr_en;

// LPD_LIN0RX interface
input             io_LPD_LIN0RX_txd;
output            io_LPD_LIN0RX_rxd;
input             io_LPD_LIN0RX_tr_en;

// EPWM0 interface
output            io_EPWM0_a_i;
input             io_EPWM0_a_o;
input             io_EPWM0_a_oen;
output            io_EPWM0_b_i;
input             io_EPWM0_b_o;
input             io_EPWM0_b_oen;

// EPWM1 interface
output            io_EPWM1_a_i;
input             io_EPWM1_a_o;
input             io_EPWM1_a_oen;
output            io_EPWM1_b_i;
input             io_EPWM1_b_o;
input             io_EPWM1_b_oen;

// EPWM2 interface
output            io_EPWM2_a_i;
input             io_EPWM2_a_o;
input             io_EPWM2_a_oen;
output            io_EPWM2_b_i;
input             io_EPWM2_b_o;
input             io_EPWM2_b_oen;

// EPWM3 interface
output            io_EPWM3_a_i;
input             io_EPWM3_a_o;
input             io_EPWM3_a_oen;
output            io_EPWM3_b_i;
input             io_EPWM3_b_o;
input             io_EPWM3_b_oen;

// EPWM4 interface
output            io_EPWM4_a_i;
input             io_EPWM4_a_o;
input             io_EPWM4_a_oen;
output            io_EPWM4_b_i;
input             io_EPWM4_b_o;
input             io_EPWM4_b_oen;

// EPWM5 interface
output            io_EPWM5_a_i;
input             io_EPWM5_a_o;
input             io_EPWM5_a_oen;
output            io_EPWM5_b_i;
input             io_EPWM5_b_o;
input             io_EPWM5_b_oen;

// EPWM6 interface
output            io_EPWM6_a_i;
input             io_EPWM6_a_o;
input             io_EPWM6_a_oen;
output            io_EPWM6_b_i;
input             io_EPWM6_b_o;
input             io_EPWM6_b_oen;

// EPWM7 interface
output            io_EPWM7_a_i;
input             io_EPWM7_a_o;
input             io_EPWM7_a_oen;
output            io_EPWM7_b_i;
input             io_EPWM7_b_o;
input             io_EPWM7_b_oen;

// EPWM8 interface
output            io_EPWM8_a_i;
input             io_EPWM8_a_o;
input             io_EPWM8_a_oen;
output            io_EPWM8_b_i;
input             io_EPWM8_b_o;
input             io_EPWM8_b_oen;

// EPWM9 interface
output            io_EPWM9_a_i;
input             io_EPWM9_a_o;
input             io_EPWM9_a_oen;
output            io_EPWM9_b_i;
input             io_EPWM9_b_o;
input             io_EPWM9_b_oen;

// EPWM10 interface
output            io_EPWM10_a_i;
input             io_EPWM10_a_o;
input             io_EPWM10_a_oen;
output            io_EPWM10_b_i;
input             io_EPWM10_b_o;
input             io_EPWM10_b_oen;

// EPWM11 interface
output            io_EPWM11_a_i;
input             io_EPWM11_a_o;
input             io_EPWM11_a_oen;
output            io_EPWM11_b_i;
input             io_EPWM11_b_o;
input             io_EPWM11_b_oen;

// EPWM12 interface
output            io_EPWM12_a_i;
input             io_EPWM12_a_o;
input             io_EPWM12_a_oen;
output            io_EPWM12_b_i;
input             io_EPWM12_b_o;
input             io_EPWM12_b_oen;

// EPWM13 interface
output            io_EPWM13_a_i;
input             io_EPWM13_a_o;
input             io_EPWM13_a_oen;
output            io_EPWM13_b_i;
input             io_EPWM13_b_o;
input             io_EPWM13_b_oen;

// EPWM14 interface
output            io_EPWM14_a_i;
input             io_EPWM14_a_o;
input             io_EPWM14_a_oen;
output            io_EPWM14_b_i;
input             io_EPWM14_b_o;
input             io_EPWM14_b_oen;

// EPWM15 interface
output            io_EPWM15_a_i;
input             io_EPWM15_a_o;
input             io_EPWM15_a_oen;
output            io_EPWM15_b_i;
input             io_EPWM15_b_o;
input             io_EPWM15_b_oen;

// EPWM16 interface
output            io_EPWM16_a_i;
input             io_EPWM16_a_o;
input             io_EPWM16_a_oen;
output            io_EPWM16_b_i;
input             io_EPWM16_b_o;
input             io_EPWM16_b_oen;

// EPWM17 interface
output            io_EPWM17_a_i;
input             io_EPWM17_a_o;
input             io_EPWM17_a_oen;
output            io_EPWM17_b_i;
input             io_EPWM17_b_o;
input             io_EPWM17_b_oen;

// EPWM18 interface
output            io_EPWM18_a_i;
input             io_EPWM18_a_o;
input             io_EPWM18_a_oen;
output            io_EPWM18_b_i;
input             io_EPWM18_b_o;
input             io_EPWM18_b_oen;

// EPWM19 interface
output            io_EPWM19_a_i;
input             io_EPWM19_a_o;
input             io_EPWM19_a_oen;
output            io_EPWM19_b_i;
input             io_EPWM19_b_o;
input             io_EPWM19_b_oen;

// EPWM20 interface
output            io_EPWM20_a_i;
input             io_EPWM20_a_o;
input             io_EPWM20_a_oen;
output            io_EPWM20_b_i;
input             io_EPWM20_b_o;
input             io_EPWM20_b_oen;

// EPWM21 interface
output            io_EPWM21_a_i;
input             io_EPWM21_a_o;
input             io_EPWM21_a_oen;
output            io_EPWM21_b_i;
input             io_EPWM21_b_o;
input             io_EPWM21_b_oen;

// EPWM22 interface
output            io_EPWM22_a_i;
input             io_EPWM22_a_o;
input             io_EPWM22_a_oen;
output            io_EPWM22_b_i;
input             io_EPWM22_b_o;
input             io_EPWM22_b_oen;

// EPWM23 interface
output            io_EPWM23_a_i;
input             io_EPWM23_a_o;
input             io_EPWM23_a_oen;
output            io_EPWM23_b_i;
input             io_EPWM23_b_o;
input             io_EPWM23_b_oen;

// EPWM24 interface
output            io_EPWM24_a_i;
input             io_EPWM24_a_o;
input             io_EPWM24_a_oen;
output            io_EPWM24_b_i;
input             io_EPWM24_b_o;
input             io_EPWM24_b_oen;

// EPWM25 interface
output            io_EPWM25_a_i;
input             io_EPWM25_a_o;
input             io_EPWM25_a_oen;
output            io_EPWM25_b_i;
input             io_EPWM25_b_o;
input             io_EPWM25_b_oen;

// EPWM26 interface
output            io_EPWM26_a_i;
input             io_EPWM26_a_o;
input             io_EPWM26_a_oen;
output            io_EPWM26_b_i;
input             io_EPWM26_b_o;
input             io_EPWM26_b_oen;

// EPWM27 interface
output            io_EPWM27_a_i;
input             io_EPWM27_a_o;
input             io_EPWM27_a_oen;
output            io_EPWM27_b_i;
input             io_EPWM27_b_o;
input             io_EPWM27_b_oen;

// EPWM28 interface
output            io_EPWM28_a_i;
input             io_EPWM28_a_o;
input             io_EPWM28_a_oen;
output            io_EPWM28_b_i;
input             io_EPWM28_b_o;
input             io_EPWM28_b_oen;

// EPWM29 interface
output            io_EPWM29_a_i;
input             io_EPWM29_a_o;
input             io_EPWM29_a_oen;
output            io_EPWM29_b_i;
input             io_EPWM29_b_o;
input             io_EPWM29_b_oen;

// EPWM30 interface
output            io_EPWM30_a_i;
input             io_EPWM30_a_o;
input             io_EPWM30_a_oen;
output            io_EPWM30_b_i;
input             io_EPWM30_b_o;
input             io_EPWM30_b_oen;

// EPWM31 interface
output            io_EPWM31_a_i;
input             io_EPWM31_a_o;
input             io_EPWM31_a_oen;
output            io_EPWM31_b_i;
input             io_EPWM31_b_o;
input             io_EPWM31_b_oen;

// EPWMSYNCO interface
output            io_EPWMSYNCO_a_i;
input             io_EPWMSYNCO_a_o;
input             io_EPWMSYNCO_a_oen;
output            io_EPWMSYNCO_b_i;
input             io_EPWMSYNCO_b_o;
input             io_EPWMSYNCO_b_oen;

// ICL  PORT
input             io_OUTPUTXBAR0_intr;

// ICL  PORT
input             io_OUTPUTXBAR1_intr;

// ICL  PORT
input             io_OUTPUTXBAR2_intr;

// ICL  PORT
input             io_OUTPUTXBAR3_intr;

// ICL  PORT
input             io_OUTPUTXBAR4_intr;

// ICL  PORT
input             io_OUTPUTXBAR5_intr;

// ICL  PORT
input             io_OUTPUTXBAR6_intr;

// ICL  PORT
input             io_OUTPUTXBAR7_intr;

// ICL  PORT
input             io_OUTPUTXBAR8_intr;

// ICL  PORT
input             io_OUTPUTXBAR9_intr;

// ICL  PORT
input             io_OUTPUTXBAR10_intr;

// ICL  PORT
input             io_OUTPUTXBAR11_intr;

// ICL  PORT
input             io_OUTPUTXBAR12_intr;

// ICL  PORT
input             io_OUTPUTXBAR13_intr;

// ICL  PORT
input             io_OUTPUTXBAR14_intr;

// ICL  PORT
input             io_OUTPUTXBAR15_intr;

// SDFM_SDFM0 interface
output            io_SDFM0_i_datain1;
output            io_SDFM0_i_clock1;
output            io_SDFM0_i_datain2;
output            io_SDFM0_i_clock2;
output            io_SDFM0_i_datain3;
output            io_SDFM0_i_clock3;
output            io_SDFM0_i_datain4;
output            io_SDFM0_i_clock4;

// SDFM_SDFM1 interface
output            io_SDFM1_i_datain1;
output            io_SDFM1_i_clock1;
output            io_SDFM1_i_datain2;
output            io_SDFM1_i_clock2;
output            io_SDFM1_i_datain3;
output            io_SDFM1_i_clock3;
output            io_SDFM1_i_datain4;
output            io_SDFM1_i_clock4;

// SDFM_SDFM2 interface
output            io_SDFM2_i_datain1;
output            io_SDFM2_i_clock1;
output            io_SDFM2_i_datain2;
output            io_SDFM2_i_clock2;
output            io_SDFM2_i_datain3;
output            io_SDFM2_i_clock3;
output            io_SDFM2_i_datain4;
output            io_SDFM2_i_clock4;

// SDFM_SDFM3 interface
output            io_SDFM3_i_datain1;
output            io_SDFM3_i_clock1;
output            io_SDFM3_i_datain2;
output            io_SDFM3_i_clock2;
output            io_SDFM3_i_datain3;
output            io_SDFM3_i_clock3;
output            io_SDFM3_i_datain4;
output            io_SDFM3_i_clock4;

// SDFM_SDFM4 interface
output            io_SDFM4_i_datain1;
output            io_SDFM4_i_clock1;
output            io_SDFM4_i_datain2;
output            io_SDFM4_i_clock2;
output            io_SDFM4_i_datain3;
output            io_SDFM4_i_clock3;
output            io_SDFM4_i_datain4;
output            io_SDFM4_i_clock4;

// SDFM_SDFM5 interface
output            io_SDFM5_i_datain1;
output            io_SDFM5_i_clock1;
output            io_SDFM5_i_datain2;
output            io_SDFM5_i_clock2;
output            io_SDFM5_i_datain3;
output            io_SDFM5_i_clock3;
output            io_SDFM5_i_datain4;
output            io_SDFM5_i_clock4;

// SDFM_SDFM6 interface
output            io_SDFM6_i_datain1;
output            io_SDFM6_i_clock1;
output            io_SDFM6_i_datain2;
output            io_SDFM6_i_clock2;
output            io_SDFM6_i_datain3;
output            io_SDFM6_i_clock3;
output            io_SDFM6_i_datain4;
output            io_SDFM6_i_clock4;

// SDFM_SDFM7 interface
output            io_SDFM7_i_datain1;
output            io_SDFM7_i_clock1;
output            io_SDFM7_i_datain2;
output            io_SDFM7_i_clock2;
output            io_SDFM7_i_datain3;
output            io_SDFM7_i_clock3;
output            io_SDFM7_i_datain4;
output            io_SDFM7_i_clock4;

// SDFM_SDFM8 interface
output            io_SDFM8_i_datain1;
output            io_SDFM8_i_clock1;
output            io_SDFM8_i_datain2;
output            io_SDFM8_i_clock2;
output            io_SDFM8_i_datain3;
output            io_SDFM8_i_clock3;
output            io_SDFM8_i_datain4;
output            io_SDFM8_i_clock4;

// SDFM_SDFM9 interface
output            io_SDFM9_i_datain1;
output            io_SDFM9_i_clock1;
output            io_SDFM9_i_datain2;
output            io_SDFM9_i_clock2;
output            io_SDFM9_i_datain3;
output            io_SDFM9_i_clock3;
output            io_SDFM9_i_datain4;
output            io_SDFM9_i_clock4;

// SDFM_SDFM10 interface
output            io_SDFM10_i_datain1;
output            io_SDFM10_i_clock1;
output            io_SDFM10_i_datain2;
output            io_SDFM10_i_clock2;
output            io_SDFM10_i_datain3;
output            io_SDFM10_i_clock3;
output            io_SDFM10_i_datain4;
output            io_SDFM10_i_clock4;

// SDFM_SDFM11 interface
output            io_SDFM11_i_datain1;
output            io_SDFM11_i_clock1;
output            io_SDFM11_i_datain2;
output            io_SDFM11_i_clock2;
output            io_SDFM11_i_datain3;
output            io_SDFM11_i_clock3;
output            io_SDFM11_i_datain4;
output            io_SDFM11_i_clock4;

// ADC0EXTMUXSEL0 interface
input       [31:0] io_ADC0EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC0EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC0EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC0EXTMUXSEL0_adcresult;
input             io_ADC0EXTMUXSEL0_adcclk;
input             io_ADC0EXTMUXSEL0_adcresolution;
input             io_ADC0EXTMUXSEL0_adcsignalmode;
input             io_ADC0EXTMUXSEL0_adcsoc;
input             io_ADC0EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC0EXTMUXSEL0_adcchsel;
input             io_ADC0EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC0EXTMUXSEL0_adccalibstep;
input             io_ADC0EXTMUXSEL0_samcapreset_disable;
input             io_ADC0EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC0EXTMUXSEL0_dtb;

// ext_ADC0EXTMUXSEL0 interface
input        [4:0] io_ext_ADC0EXTMUXSEL0_adcchsel;

// ADC0EXTMUXSEL1 interface
input       [31:0] io_ADC0EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC0EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC0EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC0EXTMUXSEL1_adcresult;
input             io_ADC0EXTMUXSEL1_adcclk;
input             io_ADC0EXTMUXSEL1_adcresolution;
input             io_ADC0EXTMUXSEL1_adcsignalmode;
input             io_ADC0EXTMUXSEL1_adcsoc;
input             io_ADC0EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC0EXTMUXSEL1_adcchsel;
input             io_ADC0EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC0EXTMUXSEL1_adccalibstep;
input             io_ADC0EXTMUXSEL1_samcapreset_disable;
input             io_ADC0EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC0EXTMUXSEL1_dtb;

// ext_ADC0EXTMUXSEL1 interface
input        [4:0] io_ext_ADC0EXTMUXSEL1_adcchsel;

// ADC0EXTMUXSEL2 interface
input       [31:0] io_ADC0EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC0EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC0EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC0EXTMUXSEL2_adcresult;
input             io_ADC0EXTMUXSEL2_adcclk;
input             io_ADC0EXTMUXSEL2_adcresolution;
input             io_ADC0EXTMUXSEL2_adcsignalmode;
input             io_ADC0EXTMUXSEL2_adcsoc;
input             io_ADC0EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC0EXTMUXSEL2_adcchsel;
input             io_ADC0EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC0EXTMUXSEL2_adccalibstep;
input             io_ADC0EXTMUXSEL2_samcapreset_disable;
input             io_ADC0EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC0EXTMUXSEL2_dtb;

// ext_ADC0EXTMUXSEL2 interface
input        [4:0] io_ext_ADC0EXTMUXSEL2_adcchsel;

// ADC0EXTMUXSEL3 interface
input       [31:0] io_ADC0EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC0EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC0EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC0EXTMUXSEL3_adcresult;
input             io_ADC0EXTMUXSEL3_adcclk;
input             io_ADC0EXTMUXSEL3_adcresolution;
input             io_ADC0EXTMUXSEL3_adcsignalmode;
input             io_ADC0EXTMUXSEL3_adcsoc;
input             io_ADC0EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC0EXTMUXSEL3_adcchsel;
input             io_ADC0EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC0EXTMUXSEL3_adccalibstep;
input             io_ADC0EXTMUXSEL3_samcapreset_disable;
input             io_ADC0EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC0EXTMUXSEL3_dtb;

// ext_ADC0EXTMUXSEL3 interface
input        [4:0] io_ext_ADC0EXTMUXSEL3_adcchsel;

// ADC1EXTMUXSEL0 interface
input       [31:0] io_ADC1EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC1EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC1EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC1EXTMUXSEL0_adcresult;
input             io_ADC1EXTMUXSEL0_adcclk;
input             io_ADC1EXTMUXSEL0_adcresolution;
input             io_ADC1EXTMUXSEL0_adcsignalmode;
input             io_ADC1EXTMUXSEL0_adcsoc;
input             io_ADC1EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC1EXTMUXSEL0_adcchsel;
input             io_ADC1EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC1EXTMUXSEL0_adccalibstep;
input             io_ADC1EXTMUXSEL0_samcapreset_disable;
input             io_ADC1EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC1EXTMUXSEL0_dtb;

// ext_ADC1EXTMUXSEL0 interface
input        [4:0] io_ext_ADC1EXTMUXSEL0_adcchsel;

// ADC1EXTMUXSEL1 interface
input       [31:0] io_ADC1EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC1EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC1EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC1EXTMUXSEL1_adcresult;
input             io_ADC1EXTMUXSEL1_adcclk;
input             io_ADC1EXTMUXSEL1_adcresolution;
input             io_ADC1EXTMUXSEL1_adcsignalmode;
input             io_ADC1EXTMUXSEL1_adcsoc;
input             io_ADC1EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC1EXTMUXSEL1_adcchsel;
input             io_ADC1EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC1EXTMUXSEL1_adccalibstep;
input             io_ADC1EXTMUXSEL1_samcapreset_disable;
input             io_ADC1EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC1EXTMUXSEL1_dtb;

// ext_ADC1EXTMUXSEL1 interface
input        [4:0] io_ext_ADC1EXTMUXSEL1_adcchsel;

// ADC1EXTMUXSEL2 interface
input       [31:0] io_ADC1EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC1EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC1EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC1EXTMUXSEL2_adcresult;
input             io_ADC1EXTMUXSEL2_adcclk;
input             io_ADC1EXTMUXSEL2_adcresolution;
input             io_ADC1EXTMUXSEL2_adcsignalmode;
input             io_ADC1EXTMUXSEL2_adcsoc;
input             io_ADC1EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC1EXTMUXSEL2_adcchsel;
input             io_ADC1EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC1EXTMUXSEL2_adccalibstep;
input             io_ADC1EXTMUXSEL2_samcapreset_disable;
input             io_ADC1EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC1EXTMUXSEL2_dtb;

// ext_ADC1EXTMUXSEL2 interface
input        [4:0] io_ext_ADC1EXTMUXSEL2_adcchsel;

// ADC1EXTMUXSEL3 interface
input       [31:0] io_ADC1EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC1EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC1EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC1EXTMUXSEL3_adcresult;
input             io_ADC1EXTMUXSEL3_adcclk;
input             io_ADC1EXTMUXSEL3_adcresolution;
input             io_ADC1EXTMUXSEL3_adcsignalmode;
input             io_ADC1EXTMUXSEL3_adcsoc;
input             io_ADC1EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC1EXTMUXSEL3_adcchsel;
input             io_ADC1EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC1EXTMUXSEL3_adccalibstep;
input             io_ADC1EXTMUXSEL3_samcapreset_disable;
input             io_ADC1EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC1EXTMUXSEL3_dtb;

// ext_ADC1EXTMUXSEL3 interface
input        [4:0] io_ext_ADC1EXTMUXSEL3_adcchsel;

// ADC2EXTMUXSEL0 interface
input       [31:0] io_ADC2EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC2EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC2EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC2EXTMUXSEL0_adcresult;
input             io_ADC2EXTMUXSEL0_adcclk;
input             io_ADC2EXTMUXSEL0_adcresolution;
input             io_ADC2EXTMUXSEL0_adcsignalmode;
input             io_ADC2EXTMUXSEL0_adcsoc;
input             io_ADC2EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC2EXTMUXSEL0_adcchsel;
input             io_ADC2EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC2EXTMUXSEL0_adccalibstep;
input             io_ADC2EXTMUXSEL0_samcapreset_disable;
input             io_ADC2EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC2EXTMUXSEL0_dtb;

// ext_ADC2EXTMUXSEL0 interface
input        [4:0] io_ext_ADC2EXTMUXSEL0_adcchsel;

// ADC2EXTMUXSEL1 interface
input       [31:0] io_ADC2EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC2EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC2EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC2EXTMUXSEL1_adcresult;
input             io_ADC2EXTMUXSEL1_adcclk;
input             io_ADC2EXTMUXSEL1_adcresolution;
input             io_ADC2EXTMUXSEL1_adcsignalmode;
input             io_ADC2EXTMUXSEL1_adcsoc;
input             io_ADC2EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC2EXTMUXSEL1_adcchsel;
input             io_ADC2EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC2EXTMUXSEL1_adccalibstep;
input             io_ADC2EXTMUXSEL1_samcapreset_disable;
input             io_ADC2EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC2EXTMUXSEL1_dtb;

// ext_ADC2EXTMUXSEL1 interface
input        [4:0] io_ext_ADC2EXTMUXSEL1_adcchsel;

// ADC2EXTMUXSEL2 interface
input       [31:0] io_ADC2EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC2EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC2EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC2EXTMUXSEL2_adcresult;
input             io_ADC2EXTMUXSEL2_adcclk;
input             io_ADC2EXTMUXSEL2_adcresolution;
input             io_ADC2EXTMUXSEL2_adcsignalmode;
input             io_ADC2EXTMUXSEL2_adcsoc;
input             io_ADC2EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC2EXTMUXSEL2_adcchsel;
input             io_ADC2EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC2EXTMUXSEL2_adccalibstep;
input             io_ADC2EXTMUXSEL2_samcapreset_disable;
input             io_ADC2EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC2EXTMUXSEL2_dtb;

// ext_ADC2EXTMUXSEL2 interface
input        [4:0] io_ext_ADC2EXTMUXSEL2_adcchsel;

// ADC2EXTMUXSEL3 interface
input       [31:0] io_ADC2EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC2EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC2EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC2EXTMUXSEL3_adcresult;
input             io_ADC2EXTMUXSEL3_adcclk;
input             io_ADC2EXTMUXSEL3_adcresolution;
input             io_ADC2EXTMUXSEL3_adcsignalmode;
input             io_ADC2EXTMUXSEL3_adcsoc;
input             io_ADC2EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC2EXTMUXSEL3_adcchsel;
input             io_ADC2EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC2EXTMUXSEL3_adccalibstep;
input             io_ADC2EXTMUXSEL3_samcapreset_disable;
input             io_ADC2EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC2EXTMUXSEL3_dtb;

// ext_ADC2EXTMUXSEL3 interface
input        [4:0] io_ext_ADC2EXTMUXSEL3_adcchsel;

// ADC3EXTMUXSEL0 interface
input       [31:0] io_ADC3EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC3EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC3EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC3EXTMUXSEL0_adcresult;
input             io_ADC3EXTMUXSEL0_adcclk;
input             io_ADC3EXTMUXSEL0_adcresolution;
input             io_ADC3EXTMUXSEL0_adcsignalmode;
input             io_ADC3EXTMUXSEL0_adcsoc;
input             io_ADC3EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC3EXTMUXSEL0_adcchsel;
input             io_ADC3EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC3EXTMUXSEL0_adccalibstep;
input             io_ADC3EXTMUXSEL0_samcapreset_disable;
input             io_ADC3EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC3EXTMUXSEL0_dtb;

// ext_ADC3EXTMUXSEL0 interface
input        [4:0] io_ext_ADC3EXTMUXSEL0_adcchsel;

// ADC3EXTMUXSEL1 interface
input       [31:0] io_ADC3EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC3EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC3EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC3EXTMUXSEL1_adcresult;
input             io_ADC3EXTMUXSEL1_adcclk;
input             io_ADC3EXTMUXSEL1_adcresolution;
input             io_ADC3EXTMUXSEL1_adcsignalmode;
input             io_ADC3EXTMUXSEL1_adcsoc;
input             io_ADC3EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC3EXTMUXSEL1_adcchsel;
input             io_ADC3EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC3EXTMUXSEL1_adccalibstep;
input             io_ADC3EXTMUXSEL1_samcapreset_disable;
input             io_ADC3EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC3EXTMUXSEL1_dtb;

// ext_ADC3EXTMUXSEL1 interface
input        [4:0] io_ext_ADC3EXTMUXSEL1_adcchsel;

// ADC3EXTMUXSEL2 interface
input       [31:0] io_ADC3EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC3EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC3EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC3EXTMUXSEL2_adcresult;
input             io_ADC3EXTMUXSEL2_adcclk;
input             io_ADC3EXTMUXSEL2_adcresolution;
input             io_ADC3EXTMUXSEL2_adcsignalmode;
input             io_ADC3EXTMUXSEL2_adcsoc;
input             io_ADC3EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC3EXTMUXSEL2_adcchsel;
input             io_ADC3EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC3EXTMUXSEL2_adccalibstep;
input             io_ADC3EXTMUXSEL2_samcapreset_disable;
input             io_ADC3EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC3EXTMUXSEL2_dtb;

// ext_ADC3EXTMUXSEL2 interface
input        [4:0] io_ext_ADC3EXTMUXSEL2_adcchsel;

// ADC3EXTMUXSEL3 interface
input       [31:0] io_ADC3EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC3EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC3EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC3EXTMUXSEL3_adcresult;
input             io_ADC3EXTMUXSEL3_adcclk;
input             io_ADC3EXTMUXSEL3_adcresolution;
input             io_ADC3EXTMUXSEL3_adcsignalmode;
input             io_ADC3EXTMUXSEL3_adcsoc;
input             io_ADC3EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC3EXTMUXSEL3_adcchsel;
input             io_ADC3EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC3EXTMUXSEL3_adccalibstep;
input             io_ADC3EXTMUXSEL3_samcapreset_disable;
input             io_ADC3EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC3EXTMUXSEL3_dtb;

// ext_ADC3EXTMUXSEL3 interface
input        [4:0] io_ext_ADC3EXTMUXSEL3_adcchsel;

// ADC4EXTMUXSEL0 interface
input       [31:0] io_ADC4EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC4EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC4EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC4EXTMUXSEL0_adcresult;
input             io_ADC4EXTMUXSEL0_adcclk;
input             io_ADC4EXTMUXSEL0_adcresolution;
input             io_ADC4EXTMUXSEL0_adcsignalmode;
input             io_ADC4EXTMUXSEL0_adcsoc;
input             io_ADC4EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC4EXTMUXSEL0_adcchsel;
input             io_ADC4EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC4EXTMUXSEL0_adccalibstep;
input             io_ADC4EXTMUXSEL0_samcapreset_disable;
input             io_ADC4EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC4EXTMUXSEL0_dtb;

// ext_ADC4EXTMUXSEL0 interface
input        [4:0] io_ext_ADC4EXTMUXSEL0_adcchsel;

// ADC4EXTMUXSEL1 interface
input       [31:0] io_ADC4EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC4EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC4EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC4EXTMUXSEL1_adcresult;
input             io_ADC4EXTMUXSEL1_adcclk;
input             io_ADC4EXTMUXSEL1_adcresolution;
input             io_ADC4EXTMUXSEL1_adcsignalmode;
input             io_ADC4EXTMUXSEL1_adcsoc;
input             io_ADC4EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC4EXTMUXSEL1_adcchsel;
input             io_ADC4EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC4EXTMUXSEL1_adccalibstep;
input             io_ADC4EXTMUXSEL1_samcapreset_disable;
input             io_ADC4EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC4EXTMUXSEL1_dtb;

// ext_ADC4EXTMUXSEL1 interface
input        [4:0] io_ext_ADC4EXTMUXSEL1_adcchsel;

// ADC4EXTMUXSEL2 interface
input       [31:0] io_ADC4EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC4EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC4EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC4EXTMUXSEL2_adcresult;
input             io_ADC4EXTMUXSEL2_adcclk;
input             io_ADC4EXTMUXSEL2_adcresolution;
input             io_ADC4EXTMUXSEL2_adcsignalmode;
input             io_ADC4EXTMUXSEL2_adcsoc;
input             io_ADC4EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC4EXTMUXSEL2_adcchsel;
input             io_ADC4EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC4EXTMUXSEL2_adccalibstep;
input             io_ADC4EXTMUXSEL2_samcapreset_disable;
input             io_ADC4EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC4EXTMUXSEL2_dtb;

// ext_ADC4EXTMUXSEL2 interface
input        [4:0] io_ext_ADC4EXTMUXSEL2_adcchsel;

// ADC4EXTMUXSEL3 interface
input       [31:0] io_ADC4EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC4EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC4EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC4EXTMUXSEL3_adcresult;
input             io_ADC4EXTMUXSEL3_adcclk;
input             io_ADC4EXTMUXSEL3_adcresolution;
input             io_ADC4EXTMUXSEL3_adcsignalmode;
input             io_ADC4EXTMUXSEL3_adcsoc;
input             io_ADC4EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC4EXTMUXSEL3_adcchsel;
input             io_ADC4EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC4EXTMUXSEL3_adccalibstep;
input             io_ADC4EXTMUXSEL3_samcapreset_disable;
input             io_ADC4EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC4EXTMUXSEL3_dtb;

// ext_ADC4EXTMUXSEL3 interface
input        [4:0] io_ext_ADC4EXTMUXSEL3_adcchsel;

// ADC5EXTMUXSEL0 interface
input       [31:0] io_ADC5EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC5EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC5EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC5EXTMUXSEL0_adcresult;
input             io_ADC5EXTMUXSEL0_adcclk;
input             io_ADC5EXTMUXSEL0_adcresolution;
input             io_ADC5EXTMUXSEL0_adcsignalmode;
input             io_ADC5EXTMUXSEL0_adcsoc;
input             io_ADC5EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC5EXTMUXSEL0_adcchsel;
input             io_ADC5EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC5EXTMUXSEL0_adccalibstep;
input             io_ADC5EXTMUXSEL0_samcapreset_disable;
input             io_ADC5EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC5EXTMUXSEL0_dtb;

// ext_ADC5EXTMUXSEL0 interface
input        [4:0] io_ext_ADC5EXTMUXSEL0_adcchsel;

// ADC5EXTMUXSEL1 interface
input       [31:0] io_ADC5EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC5EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC5EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC5EXTMUXSEL1_adcresult;
input             io_ADC5EXTMUXSEL1_adcclk;
input             io_ADC5EXTMUXSEL1_adcresolution;
input             io_ADC5EXTMUXSEL1_adcsignalmode;
input             io_ADC5EXTMUXSEL1_adcsoc;
input             io_ADC5EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC5EXTMUXSEL1_adcchsel;
input             io_ADC5EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC5EXTMUXSEL1_adccalibstep;
input             io_ADC5EXTMUXSEL1_samcapreset_disable;
input             io_ADC5EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC5EXTMUXSEL1_dtb;

// ext_ADC5EXTMUXSEL1 interface
input        [4:0] io_ext_ADC5EXTMUXSEL1_adcchsel;

// ADC5EXTMUXSEL2 interface
input       [31:0] io_ADC5EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC5EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC5EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC5EXTMUXSEL2_adcresult;
input             io_ADC5EXTMUXSEL2_adcclk;
input             io_ADC5EXTMUXSEL2_adcresolution;
input             io_ADC5EXTMUXSEL2_adcsignalmode;
input             io_ADC5EXTMUXSEL2_adcsoc;
input             io_ADC5EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC5EXTMUXSEL2_adcchsel;
input             io_ADC5EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC5EXTMUXSEL2_adccalibstep;
input             io_ADC5EXTMUXSEL2_samcapreset_disable;
input             io_ADC5EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC5EXTMUXSEL2_dtb;

// ext_ADC5EXTMUXSEL2 interface
input        [4:0] io_ext_ADC5EXTMUXSEL2_adcchsel;

// ADC5EXTMUXSEL3 interface
input       [31:0] io_ADC5EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC5EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC5EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC5EXTMUXSEL3_adcresult;
input             io_ADC5EXTMUXSEL3_adcclk;
input             io_ADC5EXTMUXSEL3_adcresolution;
input             io_ADC5EXTMUXSEL3_adcsignalmode;
input             io_ADC5EXTMUXSEL3_adcsoc;
input             io_ADC5EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC5EXTMUXSEL3_adcchsel;
input             io_ADC5EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC5EXTMUXSEL3_adccalibstep;
input             io_ADC5EXTMUXSEL3_samcapreset_disable;
input             io_ADC5EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC5EXTMUXSEL3_dtb;

// ext_ADC5EXTMUXSEL3 interface
input        [4:0] io_ext_ADC5EXTMUXSEL3_adcchsel;

// ADC6EXTMUXSEL0 interface
input       [31:0] io_ADC6EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC6EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC6EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC6EXTMUXSEL0_adcresult;
input             io_ADC6EXTMUXSEL0_adcclk;
input             io_ADC6EXTMUXSEL0_adcresolution;
input             io_ADC6EXTMUXSEL0_adcsignalmode;
input             io_ADC6EXTMUXSEL0_adcsoc;
input             io_ADC6EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC6EXTMUXSEL0_adcchsel;
input             io_ADC6EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC6EXTMUXSEL0_adccalibstep;
input             io_ADC6EXTMUXSEL0_samcapreset_disable;
input             io_ADC6EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC6EXTMUXSEL0_dtb;

// ext_ADC6EXTMUXSEL0 interface
input        [4:0] io_ext_ADC6EXTMUXSEL0_adcchsel;

// ADC6EXTMUXSEL1 interface
input       [31:0] io_ADC6EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC6EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC6EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC6EXTMUXSEL1_adcresult;
input             io_ADC6EXTMUXSEL1_adcclk;
input             io_ADC6EXTMUXSEL1_adcresolution;
input             io_ADC6EXTMUXSEL1_adcsignalmode;
input             io_ADC6EXTMUXSEL1_adcsoc;
input             io_ADC6EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC6EXTMUXSEL1_adcchsel;
input             io_ADC6EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC6EXTMUXSEL1_adccalibstep;
input             io_ADC6EXTMUXSEL1_samcapreset_disable;
input             io_ADC6EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC6EXTMUXSEL1_dtb;

// ext_ADC6EXTMUXSEL1 interface
input        [4:0] io_ext_ADC6EXTMUXSEL1_adcchsel;

// ADC6EXTMUXSEL2 interface
input       [31:0] io_ADC6EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC6EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC6EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC6EXTMUXSEL2_adcresult;
input             io_ADC6EXTMUXSEL2_adcclk;
input             io_ADC6EXTMUXSEL2_adcresolution;
input             io_ADC6EXTMUXSEL2_adcsignalmode;
input             io_ADC6EXTMUXSEL2_adcsoc;
input             io_ADC6EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC6EXTMUXSEL2_adcchsel;
input             io_ADC6EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC6EXTMUXSEL2_adccalibstep;
input             io_ADC6EXTMUXSEL2_samcapreset_disable;
input             io_ADC6EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC6EXTMUXSEL2_dtb;

// ext_ADC6EXTMUXSEL2 interface
input        [4:0] io_ext_ADC6EXTMUXSEL2_adcchsel;

// ADC6EXTMUXSEL3 interface
input       [31:0] io_ADC6EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC6EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC6EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC6EXTMUXSEL3_adcresult;
input             io_ADC6EXTMUXSEL3_adcclk;
input             io_ADC6EXTMUXSEL3_adcresolution;
input             io_ADC6EXTMUXSEL3_adcsignalmode;
input             io_ADC6EXTMUXSEL3_adcsoc;
input             io_ADC6EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC6EXTMUXSEL3_adcchsel;
input             io_ADC6EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC6EXTMUXSEL3_adccalibstep;
input             io_ADC6EXTMUXSEL3_samcapreset_disable;
input             io_ADC6EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC6EXTMUXSEL3_dtb;

// ext_ADC6EXTMUXSEL3 interface
input        [4:0] io_ext_ADC6EXTMUXSEL3_adcchsel;

// ADC7EXTMUXSEL0 interface
input       [31:0] io_ADC7EXTMUXSEL0_adcconfig;
input       [31:0] io_ADC7EXTMUXSEL0_adcinltrim1;
input       [15:0] io_ADC7EXTMUXSEL0_adcofftrim;
output      [15:0] io_ADC7EXTMUXSEL0_adcresult;
input             io_ADC7EXTMUXSEL0_adcclk;
input             io_ADC7EXTMUXSEL0_adcresolution;
input             io_ADC7EXTMUXSEL0_adcsignalmode;
input             io_ADC7EXTMUXSEL0_adcsoc;
input             io_ADC7EXTMUXSEL0_adcpwrdn;
input        [4:0] io_ADC7EXTMUXSEL0_adcchsel;
input             io_ADC7EXTMUXSEL0_adccalibmode;
input        [4:0] io_ADC7EXTMUXSEL0_adccalibstep;
input             io_ADC7EXTMUXSEL0_samcapreset_disable;
input             io_ADC7EXTMUXSEL0_samcapreset_level;
output      [15:0] io_ADC7EXTMUXSEL0_dtb;

// ext_ADC7EXTMUXSEL0 interface
input        [4:0] io_ext_ADC7EXTMUXSEL0_adcchsel;

// ADC7EXTMUXSEL1 interface
input       [31:0] io_ADC7EXTMUXSEL1_adcconfig;
input       [31:0] io_ADC7EXTMUXSEL1_adcinltrim1;
input       [15:0] io_ADC7EXTMUXSEL1_adcofftrim;
output      [15:0] io_ADC7EXTMUXSEL1_adcresult;
input             io_ADC7EXTMUXSEL1_adcclk;
input             io_ADC7EXTMUXSEL1_adcresolution;
input             io_ADC7EXTMUXSEL1_adcsignalmode;
input             io_ADC7EXTMUXSEL1_adcsoc;
input             io_ADC7EXTMUXSEL1_adcpwrdn;
input        [4:0] io_ADC7EXTMUXSEL1_adcchsel;
input             io_ADC7EXTMUXSEL1_adccalibmode;
input        [4:0] io_ADC7EXTMUXSEL1_adccalibstep;
input             io_ADC7EXTMUXSEL1_samcapreset_disable;
input             io_ADC7EXTMUXSEL1_samcapreset_level;
output      [15:0] io_ADC7EXTMUXSEL1_dtb;

// ext_ADC7EXTMUXSEL1 interface
input        [4:0] io_ext_ADC7EXTMUXSEL1_adcchsel;

// ADC7EXTMUXSEL2 interface
input       [31:0] io_ADC7EXTMUXSEL2_adcconfig;
input       [31:0] io_ADC7EXTMUXSEL2_adcinltrim1;
input       [15:0] io_ADC7EXTMUXSEL2_adcofftrim;
output      [15:0] io_ADC7EXTMUXSEL2_adcresult;
input             io_ADC7EXTMUXSEL2_adcclk;
input             io_ADC7EXTMUXSEL2_adcresolution;
input             io_ADC7EXTMUXSEL2_adcsignalmode;
input             io_ADC7EXTMUXSEL2_adcsoc;
input             io_ADC7EXTMUXSEL2_adcpwrdn;
input        [4:0] io_ADC7EXTMUXSEL2_adcchsel;
input             io_ADC7EXTMUXSEL2_adccalibmode;
input        [4:0] io_ADC7EXTMUXSEL2_adccalibstep;
input             io_ADC7EXTMUXSEL2_samcapreset_disable;
input             io_ADC7EXTMUXSEL2_samcapreset_level;
output      [15:0] io_ADC7EXTMUXSEL2_dtb;

// ext_ADC7EXTMUXSEL2 interface
input        [4:0] io_ext_ADC7EXTMUXSEL2_adcchsel;

// ADC7EXTMUXSEL3 interface
input       [31:0] io_ADC7EXTMUXSEL3_adcconfig;
input       [31:0] io_ADC7EXTMUXSEL3_adcinltrim1;
input       [15:0] io_ADC7EXTMUXSEL3_adcofftrim;
output      [15:0] io_ADC7EXTMUXSEL3_adcresult;
input             io_ADC7EXTMUXSEL3_adcclk;
input             io_ADC7EXTMUXSEL3_adcresolution;
input             io_ADC7EXTMUXSEL3_adcsignalmode;
input             io_ADC7EXTMUXSEL3_adcsoc;
input             io_ADC7EXTMUXSEL3_adcpwrdn;
input        [4:0] io_ADC7EXTMUXSEL3_adcchsel;
input             io_ADC7EXTMUXSEL3_adccalibmode;
input        [4:0] io_ADC7EXTMUXSEL3_adccalibstep;
input             io_ADC7EXTMUXSEL3_samcapreset_disable;
input             io_ADC7EXTMUXSEL3_samcapreset_level;
output      [15:0] io_ADC7EXTMUXSEL3_dtb;

// ext_ADC7EXTMUXSEL3 interface
input        [4:0] io_ext_ADC7EXTMUXSEL3_adcchsel;

// ADCSOC0 interface
input       [31:0] io_ADCSOC0_adcconfig;
input       [31:0] io_ADCSOC0_adcinltrim1;
input       [15:0] io_ADCSOC0_adcofftrim;
output      [15:0] io_ADCSOC0_adcresult;
input             io_ADCSOC0_adcclk;
input             io_ADCSOC0_adcresolution;
input             io_ADCSOC0_adcsignalmode;
input             io_ADCSOC0_adcsoc;
input             io_ADCSOC0_adcpwrdn;
input        [4:0] io_ADCSOC0_adcchsel;
input             io_ADCSOC0_adccalibmode;
input        [4:0] io_ADCSOC0_adccalibstep;
input             io_ADCSOC0_samcapreset_disable;
input             io_ADCSOC0_samcapreset_level;
output      [15:0] io_ADCSOC0_dtb;

// ext_ADCSOC0 interface
input        [4:0] io_ext_ADCSOC0_adcchsel;

// ADCSOC1 interface
input       [31:0] io_ADCSOC1_adcconfig;
input       [31:0] io_ADCSOC1_adcinltrim1;
input       [15:0] io_ADCSOC1_adcofftrim;
output      [15:0] io_ADCSOC1_adcresult;
input             io_ADCSOC1_adcclk;
input             io_ADCSOC1_adcresolution;
input             io_ADCSOC1_adcsignalmode;
input             io_ADCSOC1_adcsoc;
input             io_ADCSOC1_adcpwrdn;
input        [4:0] io_ADCSOC1_adcchsel;
input             io_ADCSOC1_adccalibmode;
input        [4:0] io_ADCSOC1_adccalibstep;
input             io_ADCSOC1_samcapreset_disable;
input             io_ADCSOC1_samcapreset_level;
output      [15:0] io_ADCSOC1_dtb;

// ext_ADCSOC1 interface
input        [4:0] io_ext_ADCSOC1_adcchsel;

// FSI0TX interface
input             io_FSI0TX_ck;
input             io_FSI0TX_d0;
input             io_FSI0TX_d1;

// FSI0RX interface
output            io_FSI0RX_ck;
output            io_FSI0RX_d0;
output            io_FSI0RX_d1;

// FSI1TX interface
input             io_FSI1TX_ck;
input             io_FSI1TX_d0;
input             io_FSI1TX_d1;

// FSI1RX interface
output            io_FSI1RX_ck;
output            io_FSI1RX_d0;
output            io_FSI1RX_d1;

// FSI2TX interface
input             io_FSI2TX_ck;
input             io_FSI2TX_d0;
input             io_FSI2TX_d1;

// FSI2RX interface
output            io_FSI2RX_ck;
output            io_FSI2RX_d0;
output            io_FSI2RX_d1;

// FSI3TX interface
input             io_FSI3TX_ck;
input             io_FSI3TX_d0;
input             io_FSI3TX_d1;

// FSI3RX interface
output            io_FSI3RX_ck;
output            io_FSI3RX_d0;
output            io_FSI3RX_d1;

// FSI4TX interface
input             io_FSI4TX_ck;
input             io_FSI4TX_d0;
input             io_FSI4TX_d1;

// FSI4RX interface
output            io_FSI4RX_ck;
output            io_FSI4RX_d0;
output            io_FSI4RX_d1;

// FSI5TX interface
input             io_FSI5TX_ck;
input             io_FSI5TX_d0;
input             io_FSI5TX_d1;

// FSI5RX interface
output            io_FSI5RX_ck;
output            io_FSI5RX_d0;
output            io_FSI5RX_d1;

// I2C0SCL interface
output            io_I2C0SCL_piscl;
output            io_I2C0SCL_pisda;
input             io_I2C0SCL_porscl;
input             io_I2C0SCL_porsda;
input             io_I2C0SCL_porsccbe;
input             io_I2C0SCL_porsclhsmode;
input             io_I2C0SCL_porsclnmode;
input             io_I2C0SCL_porsdhsmode;
input             io_I2C0SCL_porsdanmode;
input             io_I2C0SCL_porsdagzn;

// I2C1SCL interface
output            io_I2C1SCL_piscl;
output            io_I2C1SCL_pisda;
input             io_I2C1SCL_porscl;
input             io_I2C1SCL_porsda;
input             io_I2C1SCL_porsccbe;
input             io_I2C1SCL_porsclhsmode;
input             io_I2C1SCL_porsclnmode;
input             io_I2C1SCL_porsdhsmode;
input             io_I2C1SCL_porsdanmode;
input             io_I2C1SCL_porsdagzn;

// I2C2SCL interface
output            io_I2C2SCL_piscl;
output            io_I2C2SCL_pisda;
input             io_I2C2SCL_porscl;
input             io_I2C2SCL_porsda;
input             io_I2C2SCL_porsccbe;
input             io_I2C2SCL_porsclhsmode;
input             io_I2C2SCL_porsclnmode;
input             io_I2C2SCL_porsdhsmode;
input             io_I2C2SCL_porsdanmode;
input             io_I2C2SCL_porsdagzn;

// I2C3SCL interface
output            io_I2C3SCL_piscl;
output            io_I2C3SCL_pisda;
input             io_I2C3SCL_porscl;
input             io_I2C3SCL_porsda;
input             io_I2C3SCL_porsccbe;
input             io_I2C3SCL_porsclhsmode;
input             io_I2C3SCL_porsclnmode;
input             io_I2C3SCL_porsdhsmode;
input             io_I2C3SCL_porsdanmode;
input             io_I2C3SCL_porsdagzn;

// XSPI0 interface
output            io_XSPI0_mst_in_clk;
input             io_XSPI0_out_clk;
input        [3:0] io_XSPI0_cs_o;
output       [7:0] io_XSPI0_data_i;
input        [7:0] io_XSPI0_data_o;
input        [7:0] io_XSPI0_data_oe_n;
input             io_XSPI0_data_mask_o;
input             io_XSPI0_data_mask_oe_n;
input        [3:0] io_XSPI0_reset_out;
output       [3:0] io_XSPI0_reset_in;
output       [3:0] io_XSPI0_intr_n;
output            io_XSPI0_dqs_clk;

// CAN0 interface
input             io_CAN0_txd;
output            io_CAN0_rxd;

// CAN1 interface
input             io_CAN1_txd;
output            io_CAN1_rxd;

// CAN2 interface
input             io_CAN2_txd;
output            io_CAN2_rxd;

// CAN3 interface
input             io_CAN3_txd;
output            io_CAN3_rxd;

// CAN4 interface
input             io_CAN4_txd;
output            io_CAN4_rxd;

// CAN5 interface
input             io_CAN5_txd;
output            io_CAN5_rxd;

// CAN6 interface
input             io_CAN6_txd;
output            io_CAN6_rxd;

// CAN7 interface
input             io_CAN7_txd;
output            io_CAN7_rxd;

// CAN8 interface
input             io_CAN8_txd;
output            io_CAN8_rxd;

// CAN9 interface
input             io_CAN9_txd;
output            io_CAN9_rxd;

// CAN10 interface
input             io_CAN10_txd;
output            io_CAN10_rxd;

// CAN11 interface
input             io_CAN11_txd;
output            io_CAN11_rxd;

// LIN0 interface
input             io_LIN0_txd;
output            io_LIN0_rxd;
input             io_LIN0_tr_en;

// LIN1 interface
input             io_LIN1_txd;
output            io_LIN1_rxd;
input             io_LIN1_tr_en;

// LIN2 interface
input             io_LIN2_txd;
output            io_LIN2_rxd;
input             io_LIN2_tr_en;

// LIN3 interface
input             io_LIN3_txd;
output            io_LIN3_rxd;
input             io_LIN3_tr_en;

// LIN4 interface
input             io_LIN4_txd;
output            io_LIN4_rxd;
input             io_LIN4_tr_en;

// LIN5 interface
input             io_LIN5_txd;
output            io_LIN5_rxd;
input             io_LIN5_tr_en;

// LIN6 interface
input             io_LIN6_txd;
output            io_LIN6_rxd;
input             io_LIN6_tr_en;

// LIN7 interface
input             io_LIN7_txd;
output            io_LIN7_rxd;
input             io_LIN7_tr_en;

// UART_IO interface
output            io_UART0_cd_n;
output            io_UART0_cts_n;
output            io_UART0_dsr_n;
input             io_UART0_dtr_n;
input             io_UART0_out1;
input             io_UART0_out2;
output            io_UART0_ri_n;
input             io_UART0_rts_n;
output            io_UART0_rx;
input             io_UART0_tx;

// UART_IO interface
output            io_UART1_cd_n;
output            io_UART1_cts_n;
output            io_UART1_dsr_n;
input             io_UART1_dtr_n;
input             io_UART1_out1;
input             io_UART1_out2;
output            io_UART1_ri_n;
input             io_UART1_rts_n;
output            io_UART1_rx;
input             io_UART1_tx;

// SENT0 interface
input      [121:0] io_SENT0_soc_ext_trig_i;
input       [31:0] io_SENT0_tstamp_val_i;
input             io_SENT0_rxd_i;
output            io_SENT0_rxd_o;
output            io_SENT0_rxd_oen_o;

// SENT1 interface
input      [121:0] io_SENT1_soc_ext_trig_i;
input       [31:0] io_SENT1_tstamp_val_i;
input             io_SENT1_rxd_i;
output            io_SENT1_rxd_o;
output            io_SENT1_rxd_oen_o;

// SENT2 interface
input      [121:0] io_SENT2_soc_ext_trig_i;
input       [31:0] io_SENT2_tstamp_val_i;
input             io_SENT2_rxd_i;
output            io_SENT2_rxd_o;
output            io_SENT2_rxd_oen_o;

// SENT3 interface
input      [121:0] io_SENT3_soc_ext_trig_i;
input       [31:0] io_SENT3_tstamp_val_i;
input             io_SENT3_rxd_i;
output            io_SENT3_rxd_o;
output            io_SENT3_rxd_oen_o;

// SENT4 interface
input      [121:0] io_SENT4_soc_ext_trig_i;
input       [31:0] io_SENT4_tstamp_val_i;
input             io_SENT4_rxd_i;
output            io_SENT4_rxd_o;
output            io_SENT4_rxd_oen_o;

// SENT5 interface
input      [121:0] io_SENT5_soc_ext_trig_i;
input       [31:0] io_SENT5_tstamp_val_i;
input             io_SENT5_rxd_i;
output            io_SENT5_rxd_o;
output            io_SENT5_rxd_oen_o;

// MIBSPI0CLK interface
input             io_MIBSPI0CLK_clock;

// MIBSPI0PICO interface
output            io_MIBSPI0PICO_in;
input             io_MIBSPI0PICO_out;
input             io_MIBSPI0PICO_oen;

// MIBSPI0POCI interface
output            io_MIBSPI0POCI_in;
input             io_MIBSPI0POCI_out;
input             io_MIBSPI0POCI_oen;

// MIBSPI0CS0 interface
output            io_MIBSPI0CS0_in;
input             io_MIBSPI0CS0_out;
input             io_MIBSPI0CS0_oen;

// MIBSPI0CS1 interface
output            io_MIBSPI0CS1_in;
input             io_MIBSPI0CS1_out;
input             io_MIBSPI0CS1_oen;

// MIBSPI0CS2 interface
output            io_MIBSPI0CS2_in;
input             io_MIBSPI0CS2_out;
input             io_MIBSPI0CS2_oen;

// MIBSPI0CS3 interface
output            io_MIBSPI0CS3_in;
input             io_MIBSPI0CS3_out;
input             io_MIBSPI0CS3_oen;

// MIBSPI0CS4 interface
output            io_MIBSPI0CS4_in;
input             io_MIBSPI0CS4_out;
input             io_MIBSPI0CS4_oen;

// MIBSPI0CS5 interface
output            io_MIBSPI0CS5_in;
input             io_MIBSPI0CS5_out;
input             io_MIBSPI0CS5_oen;

// MIBSPI0CS6 interface
output            io_MIBSPI0CS6_in;
input             io_MIBSPI0CS6_out;
input             io_MIBSPI0CS6_oen;

// MIBSPI0CS7 interface
output            io_MIBSPI0CS7_in;
input             io_MIBSPI0CS7_out;
input             io_MIBSPI0CS7_oen;

// MIBSPI0CS8 interface
output            io_MIBSPI0CS8_in;
input             io_MIBSPI0CS8_out;
input             io_MIBSPI0CS8_oen;

// MIBSPI0CS9 interface
output            io_MIBSPI0CS9_in;
input             io_MIBSPI0CS9_out;
input             io_MIBSPI0CS9_oen;

// MIBSPI0CS10 interface
output            io_MIBSPI0CS10_in;
input             io_MIBSPI0CS10_out;
input             io_MIBSPI0CS10_oen;

// MIBSPI0CS11 interface
output            io_MIBSPI0CS11_in;
input             io_MIBSPI0CS11_out;
input             io_MIBSPI0CS11_oen;

// MIBSPI1CLK interface
input             io_MIBSPI1CLK_clock;

// MIBSPI1PICO interface
output            io_MIBSPI1PICO_in;
input             io_MIBSPI1PICO_out;
input             io_MIBSPI1PICO_oen;

// MIBSPI1POCI interface
output            io_MIBSPI1POCI_in;
input             io_MIBSPI1POCI_out;
input             io_MIBSPI1POCI_oen;

// MIBSPI1CS0 interface
output            io_MIBSPI1CS0_in;
input             io_MIBSPI1CS0_out;
input             io_MIBSPI1CS0_oen;

// MIBSPI1CS1 interface
output            io_MIBSPI1CS1_in;
input             io_MIBSPI1CS1_out;
input             io_MIBSPI1CS1_oen;

// MIBSPI1CS2 interface
output            io_MIBSPI1CS2_in;
input             io_MIBSPI1CS2_out;
input             io_MIBSPI1CS2_oen;

// MIBSPI1CS3 interface
output            io_MIBSPI1CS3_in;
input             io_MIBSPI1CS3_out;
input             io_MIBSPI1CS3_oen;

// MIBSPI1CS4 interface
output            io_MIBSPI1CS4_in;
input             io_MIBSPI1CS4_out;
input             io_MIBSPI1CS4_oen;

// MIBSPI1CS5 interface
output            io_MIBSPI1CS5_in;
input             io_MIBSPI1CS5_out;
input             io_MIBSPI1CS5_oen;

// MIBSPI1CS6 interface
output            io_MIBSPI1CS6_in;
input             io_MIBSPI1CS6_out;
input             io_MIBSPI1CS6_oen;

// MIBSPI1CS7 interface
output            io_MIBSPI1CS7_in;
input             io_MIBSPI1CS7_out;
input             io_MIBSPI1CS7_oen;

// MIBSPI1CS8 interface
output            io_MIBSPI1CS8_in;
input             io_MIBSPI1CS8_out;
input             io_MIBSPI1CS8_oen;

// MIBSPI1CS9 interface
output            io_MIBSPI1CS9_in;
input             io_MIBSPI1CS9_out;
input             io_MIBSPI1CS9_oen;

// MIBSPI1CS10 interface
output            io_MIBSPI1CS10_in;
input             io_MIBSPI1CS10_out;
input             io_MIBSPI1CS10_oen;

// MIBSPI1CS11 interface
output            io_MIBSPI1CS11_in;
input             io_MIBSPI1CS11_out;
input             io_MIBSPI1CS11_oen;

// SPI2CLK interface
input             io_SPI2CLK_clock;

// SPI2PICO interface
output            io_SPI2PICO_in;
input             io_SPI2PICO_out;
input             io_SPI2PICO_oen;

// SPI2POCI interface
output            io_SPI2POCI_in;
input             io_SPI2POCI_out;
input             io_SPI2POCI_oen;

// SPI2CS0 interface
output            io_SPI2CS0_in;
input             io_SPI2CS0_out;
input             io_SPI2CS0_oen;

// SPI2CS1 interface
output            io_SPI2CS1_in;
input             io_SPI2CS1_out;
input             io_SPI2CS1_oen;

// SPI2CS2 interface
output            io_SPI2CS2_in;
input             io_SPI2CS2_out;
input             io_SPI2CS2_oen;

// SPI2CS3 interface
output            io_SPI2CS3_in;
input             io_SPI2CS3_out;
input             io_SPI2CS3_oen;

// SPI2CS4 interface
output            io_SPI2CS4_in;
input             io_SPI2CS4_out;
input             io_SPI2CS4_oen;

// SPI2CS5 interface
output            io_SPI2CS5_in;
input             io_SPI2CS5_out;
input             io_SPI2CS5_oen;

// SPI3CLK interface
input             io_SPI3CLK_clock;

// SPI3PICO interface
output            io_SPI3PICO_in;
input             io_SPI3PICO_out;
input             io_SPI3PICO_oen;

// SPI3POCI interface
output            io_SPI3POCI_in;
input             io_SPI3POCI_out;
input             io_SPI3POCI_oen;

// SPI3CS0 interface
output            io_SPI3CS0_in;
input             io_SPI3CS0_out;
input             io_SPI3CS0_oen;

// SPI3CS1 interface
output            io_SPI3CS1_in;
input             io_SPI3CS1_out;
input             io_SPI3CS1_oen;

// SPI3CS2 interface
output            io_SPI3CS2_in;
input             io_SPI3CS2_out;
input             io_SPI3CS2_oen;

// SPI3CS3 interface
output            io_SPI3CS3_in;
input             io_SPI3CS3_out;
input             io_SPI3CS3_oen;

// SPI3CS4 interface
output            io_SPI3CS4_in;
input             io_SPI3CS4_out;
input             io_SPI3CS4_oen;

// SPI3CS5 interface
output            io_SPI3CS5_in;
input             io_SPI3CS5_out;
input             io_SPI3CS5_oen;

// SPI4CLK interface
input             io_SPI4CLK_clock;

// SPI4PICO interface
output            io_SPI4PICO_in;
input             io_SPI4PICO_out;
input             io_SPI4PICO_oen;

// SPI4POCI interface
output            io_SPI4POCI_in;
input             io_SPI4POCI_out;
input             io_SPI4POCI_oen;

// SPI4CS0 interface
output            io_SPI4CS0_in;
input             io_SPI4CS0_out;
input             io_SPI4CS0_oen;

// SPI4CS1 interface
output            io_SPI4CS1_in;
input             io_SPI4CS1_out;
input             io_SPI4CS1_oen;

// SPI4CS2 interface
output            io_SPI4CS2_in;
input             io_SPI4CS2_out;
input             io_SPI4CS2_oen;

// SPI4CS3 interface
output            io_SPI4CS3_in;
input             io_SPI4CS3_out;
input             io_SPI4CS3_oen;

// SPI4CS4 interface
output            io_SPI4CS4_in;
input             io_SPI4CS4_out;
input             io_SPI4CS4_oen;

// SPI4CS5 interface
output            io_SPI4CS5_in;
input             io_SPI4CS5_out;
input             io_SPI4CS5_oen;

// SPI5CLK interface
input             io_SPI5CLK_clock;

// SPI5PICO interface
output            io_SPI5PICO_in;
input             io_SPI5PICO_out;
input             io_SPI5PICO_oen;

// SPI5POCI interface
output            io_SPI5POCI_in;
input             io_SPI5POCI_out;
input             io_SPI5POCI_oen;

// SPI5CS0 interface
output            io_SPI5CS0_in;
input             io_SPI5CS0_out;
input             io_SPI5CS0_oen;

// SPI5CS1 interface
output            io_SPI5CS1_in;
input             io_SPI5CS1_out;
input             io_SPI5CS1_oen;

// SPI5CS2 interface
output            io_SPI5CS2_in;
input             io_SPI5CS2_out;
input             io_SPI5CS2_oen;

// SPI5CS3 interface
output            io_SPI5CS3_in;
input             io_SPI5CS3_out;
input             io_SPI5CS3_oen;

// SPI5CS4 interface
output            io_SPI5CS4_in;
input             io_SPI5CS4_out;
input             io_SPI5CS4_oen;

// SPI5CS5 interface
output            io_SPI5CS5_in;
input             io_SPI5CS5_out;
input             io_SPI5CS5_oen;

// SPI6CLK interface
input             io_SPI6CLK_clock;

// SPI6PICO interface
output            io_SPI6PICO_in;
input             io_SPI6PICO_out;
input             io_SPI6PICO_oen;

// SPI6POCI interface
output            io_SPI6POCI_in;
input             io_SPI6POCI_out;
input             io_SPI6POCI_oen;

// SPI6CS0 interface
output            io_SPI6CS0_in;
input             io_SPI6CS0_out;
input             io_SPI6CS0_oen;

// SPI6CS1 interface
output            io_SPI6CS1_in;
input             io_SPI6CS1_out;
input             io_SPI6CS1_oen;

// SPI6CS2 interface
output            io_SPI6CS2_in;
input             io_SPI6CS2_out;
input             io_SPI6CS2_oen;

// SPI6CS3 interface
output            io_SPI6CS3_in;
input             io_SPI6CS3_out;
input             io_SPI6CS3_oen;

// SPI6CS4 interface
output            io_SPI6CS4_in;
input             io_SPI6CS4_out;
input             io_SPI6CS4_oen;

// SPI6CS5 interface
output            io_SPI6CS5_in;
input             io_SPI6CS5_out;
input             io_SPI6CS5_oen;

// SPI7CLK interface
input             io_SPI7CLK_clock;

// SPI7PICO interface
output            io_SPI7PICO_in;
input             io_SPI7PICO_out;
input             io_SPI7PICO_oen;

// SPI7POCI interface
output            io_SPI7POCI_in;
input             io_SPI7POCI_out;
input             io_SPI7POCI_oen;

// SPI7CS0 interface
output            io_SPI7CS0_in;
input             io_SPI7CS0_out;
input             io_SPI7CS0_oen;

// SPI7CS1 interface
output            io_SPI7CS1_in;
input             io_SPI7CS1_out;
input             io_SPI7CS1_oen;

// SPI7CS2 interface
output            io_SPI7CS2_in;
input             io_SPI7CS2_out;
input             io_SPI7CS2_oen;

// SPI7CS3 interface
output            io_SPI7CS3_in;
input             io_SPI7CS3_out;
input             io_SPI7CS3_oen;

// SPI7CS4 interface
output            io_SPI7CS4_in;
input             io_SPI7CS4_out;
input             io_SPI7CS4_oen;

// SPI7CS5 interface
output            io_SPI7CS5_in;
input             io_SPI7CS5_out;
input             io_SPI7CS5_oen;

// SPI8CLK interface
input             io_SPI8CLK_clock;

// SPI8PICO interface
output            io_SPI8PICO_in;
input             io_SPI8PICO_out;
input             io_SPI8PICO_oen;

// SPI8POCI interface
output            io_SPI8POCI_in;
input             io_SPI8POCI_out;
input             io_SPI8POCI_oen;

// SPI8CS0 interface
output            io_SPI8CS0_in;
input             io_SPI8CS0_out;
input             io_SPI8CS0_oen;

// SPI8CS1 interface
output            io_SPI8CS1_in;
input             io_SPI8CS1_out;
input             io_SPI8CS1_oen;

// SPI8CS2 interface
output            io_SPI8CS2_in;
input             io_SPI8CS2_out;
input             io_SPI8CS2_oen;

// SPI8CS3 interface
output            io_SPI8CS3_in;
input             io_SPI8CS3_out;
input             io_SPI8CS3_oen;

// SPI8CS4 interface
output            io_SPI8CS4_in;
input             io_SPI8CS4_out;
input             io_SPI8CS4_oen;

// SPI8CS5 interface
output            io_SPI8CS5_in;
input             io_SPI8CS5_out;
input             io_SPI8CS5_oen;

// SPI9CLK interface
input             io_SPI9CLK_clock;

// SPI9PICO interface
output            io_SPI9PICO_in;
input             io_SPI9PICO_out;
input             io_SPI9PICO_oen;

// SPI9POCI interface
output            io_SPI9POCI_in;
input             io_SPI9POCI_out;
input             io_SPI9POCI_oen;

// SPI9CS0 interface
output            io_SPI9CS0_in;
input             io_SPI9CS0_out;
input             io_SPI9CS0_oen;

// SPI9CS1 interface
output            io_SPI9CS1_in;
input             io_SPI9CS1_out;
input             io_SPI9CS1_oen;

// SPI9CS2 interface
output            io_SPI9CS2_in;
input             io_SPI9CS2_out;
input             io_SPI9CS2_oen;

// SPI9CS3 interface
output            io_SPI9CS3_in;
input             io_SPI9CS3_out;
input             io_SPI9CS3_oen;

// SPI9CS4 interface
output            io_SPI9CS4_in;
input             io_SPI9CS4_out;
input             io_SPI9CS4_oen;

// SPI9CS5 interface
output            io_SPI9CS5_in;
input             io_SPI9CS5_out;
input             io_SPI9CS5_oen;

// PSI5_IO interface
input        [3:0] io_PSI5_0_tx;
output       [3:0] io_PSI5_0_rx;

// PSI5_IO interface
input        [3:0] io_PSI5_1_tx;
output       [3:0] io_PSI5_1_rx;

// PSI5_IO interface
input        [3:0] io_PSI5_2_tx;
output       [3:0] io_PSI5_2_rx;

// PSI5_IO interface
input        [3:0] io_PSI5_3_tx;
output       [3:0] io_PSI5_3_rx;

//======================================
// Signal Declarations
//======================================
wire            AP0_0_IO;
wire            AP0_10_IO;
wire            AP0_11_IO;
wire            AP0_12_IO;
wire            AP0_13_IO;
wire            AP0_14_IO;
wire            AP0_15_IO;
wire            AP0_16_IO;
wire            AP0_17_IO;
wire            AP0_18_IO;
wire            AP0_19_IO;
wire            AP0_1_IO;
wire            AP0_20_IO;
wire            AP0_21_IO;
wire            AP0_22_IO;
wire            AP0_23_IO;
wire            AP0_24_IO;
wire            AP0_25_IO;
wire            AP0_26_IO;
wire            AP0_27_IO;
wire            AP0_28_IO;
wire            AP0_29_IO;
wire            AP0_2_IO;
wire            AP0_30_IO;
wire            AP0_31_IO;
wire            AP0_3_IO;
wire            AP0_4_IO;
wire            AP0_5_IO;
wire            AP0_6_IO;
wire            AP0_7_IO;
wire            AP0_8_IO;
wire            AP0_9_IO;
wire            AP0_IO;
wire            AP10_IO;
wire            AP11_IO;
wire            AP12_IO;
wire            AP13_IO;
wire            AP14_IO;
wire            AP15_IO;
wire            AP16_IO;
wire            AP17_IO;
wire            AP18_IO;
wire            AP19_IO;
wire            AP1_0_IO;
wire            AP1_10_IO;
wire            AP1_11_IO;
wire            AP1_12_IO;
wire            AP1_13_IO;
wire            AP1_14_IO;
wire            AP1_15_IO;
wire            AP1_1_IO;
wire            AP1_2_IO;
wire            AP1_3_IO;
wire            AP1_4_IO;
wire            AP1_5_IO;
wire            AP1_6_IO;
wire            AP1_7_IO;
wire            AP1_8_IO;
wire            AP1_9_IO;
wire            AP1_IO;
wire            AP20_IO;
wire            AP21_IO;
wire            AP22_IO;
wire            AP23_IO;
wire            AP24_IO;
wire            AP25_IO;
wire            AP26_IO;
wire            AP27_IO;
wire            AP28_IO;
wire            AP29_IO;
wire            AP2_IO;
wire            AP30_IO;
wire            AP31_IO;
wire            AP32_IO;
wire            AP33_IO;
wire            AP34_IO;
wire            AP35_IO;
wire            AP36_IO;
wire            AP37_IO;
wire            AP38_IO;
wire            AP39_IO;
wire            AP3_IO;
wire            AP40_IO;
wire            AP41_IO;
wire            AP42_IO;
wire            AP43_IO;
wire            AP44_IO;
wire            AP45_IO;
wire            AP46_IO;
wire            AP47_IO;
wire            AP4_IO;
wire            AP5_IO;
wire            AP6_IO;
wire            AP7_IO;
wire            AP8_IO;
wire            AP9_IO;
wire            AURORACLKN_IO;
wire            AURORACLKP_IO;
wire            AURORADN_IO;
wire            AURORADP_IO;
wire            DCDCNMOS_IO;
wire            DCDCPMOS_IO;
wire            DP0_0_IO;
wire      [7:0] DP0_0_in_mux_en_mscbus;
wire      [7:0] DP0_0_in_mux_peripheral_mscbus;
wire            DP0_0_out_demux_peripheral_mscbus;
wire            DP0_10_IO;
wire      [6:0] DP0_10_in_mux_en_mscbus;
wire      [6:0] DP0_10_in_mux_peripheral_mscbus;
wire      [1:0] DP0_10_out_demux_peripheral_mscbus;
wire            DP0_11_IO;
wire      [6:0] DP0_11_in_mux_en_mscbus;
wire      [6:0] DP0_11_in_mux_peripheral_mscbus;
wire      [1:0] DP0_11_out_demux_peripheral_mscbus;
wire            DP0_12_IO;
wire      [6:0] DP0_12_in_mux_en_mscbus;
wire      [6:0] DP0_12_in_mux_peripheral_mscbus;
wire      [1:0] DP0_12_out_demux_peripheral_mscbus;
wire            DP0_13_IO;
wire      [6:0] DP0_13_in_mux_en_mscbus;
wire      [6:0] DP0_13_in_mux_peripheral_mscbus;
wire      [2:0] DP0_13_out_demux_peripheral_mscbus;
wire            DP0_14_IO;
wire      [6:0] DP0_14_in_mux_en_mscbus;
wire      [6:0] DP0_14_in_mux_peripheral_mscbus;
wire      [1:0] DP0_14_out_demux_peripheral_mscbus;
wire            DP0_15_IO;
wire      [6:0] DP0_15_in_mux_en_mscbus;
wire      [6:0] DP0_15_in_mux_peripheral_mscbus;
wire      [1:0] DP0_15_out_demux_peripheral_mscbus;
wire            DP0_16_IO;
wire      [5:0] DP0_16_in_mux_en_mscbus;
wire      [5:0] DP0_16_in_mux_peripheral_mscbus;
wire      [3:0] DP0_16_out_demux_peripheral_mscbus;
wire            DP0_17_IO;
wire      [6:0] DP0_17_in_mux_en_mscbus;
wire      [6:0] DP0_17_in_mux_peripheral_mscbus;
wire      [2:0] DP0_17_out_demux_peripheral_mscbus;
wire            DP0_18_IO;
wire      [6:0] DP0_18_in_mux_en_mscbus;
wire      [6:0] DP0_18_in_mux_peripheral_mscbus;
wire      [2:0] DP0_18_out_demux_peripheral_mscbus;
wire            DP0_19_IO;
wire      [7:0] DP0_19_in_mux_en_mscbus;
wire      [7:0] DP0_19_in_mux_peripheral_mscbus;
wire      [1:0] DP0_19_out_demux_peripheral_mscbus;
wire            DP0_1_IO;
wire      [5:0] DP0_1_in_mux_en_mscbus;
wire      [5:0] DP0_1_in_mux_peripheral_mscbus;
wire      [3:0] DP0_1_out_demux_peripheral_mscbus;
wire            DP0_20_IO;
wire      [6:0] DP0_20_in_mux_en_mscbus;
wire      [6:0] DP0_20_in_mux_peripheral_mscbus;
wire            DP0_20_out_demux_peripheral_mscbus;
wire            DP0_21_IO;
wire      [5:0] DP0_21_in_mux_en_mscbus;
wire      [5:0] DP0_21_in_mux_peripheral_mscbus;
wire      [1:0] DP0_21_out_demux_peripheral_mscbus;
wire            DP0_22_IO;
wire      [4:0] DP0_22_in_mux_en_mscbus;
wire      [4:0] DP0_22_in_mux_peripheral_mscbus;
wire      [2:0] DP0_22_out_demux_peripheral_mscbus;
wire            DP0_23_IO;
wire      [4:0] DP0_23_in_mux_en_mscbus;
wire      [4:0] DP0_23_in_mux_peripheral_mscbus;
wire      [2:0] DP0_23_out_demux_peripheral_mscbus;
wire            DP0_24_IO;
wire      [4:0] DP0_24_in_mux_en_mscbus;
wire      [4:0] DP0_24_in_mux_peripheral_mscbus;
wire      [2:0] DP0_24_out_demux_peripheral_mscbus;
wire            DP0_25_IO;
wire      [5:0] DP0_25_in_mux_en_mscbus;
wire      [5:0] DP0_25_in_mux_peripheral_mscbus;
wire      [1:0] DP0_25_out_demux_peripheral_mscbus;
wire            DP0_26_IO;
wire      [5:0] DP0_26_in_mux_en_mscbus;
wire      [5:0] DP0_26_in_mux_peripheral_mscbus;
wire      [1:0] DP0_26_out_demux_peripheral_mscbus;
wire            DP0_27_IO;
wire      [5:0] DP0_27_in_mux_en_mscbus;
wire      [5:0] DP0_27_in_mux_peripheral_mscbus;
wire      [1:0] DP0_27_out_demux_peripheral_mscbus;
wire            DP0_28_IO;
wire      [4:0] DP0_28_in_mux_en_mscbus;
wire      [4:0] DP0_28_in_mux_peripheral_mscbus;
wire      [1:0] DP0_28_out_demux_peripheral_mscbus;
wire            DP0_29_IO;
wire      [3:0] DP0_29_in_mux_en_mscbus;
wire      [3:0] DP0_29_in_mux_peripheral_mscbus;
wire      [2:0] DP0_29_out_demux_peripheral_mscbus;
wire            DP0_2_IO;
wire      [6:0] DP0_2_in_mux_en_mscbus;
wire      [6:0] DP0_2_in_mux_peripheral_mscbus;
wire            DP0_2_out_demux_peripheral_mscbus;
wire            DP0_30_IO;
wire      [3:0] DP0_30_in_mux_en_mscbus;
wire      [3:0] DP0_30_in_mux_peripheral_mscbus;
wire      [2:0] DP0_30_out_demux_peripheral_mscbus;
wire            DP0_31_IO;
wire      [4:0] DP0_31_in_mux_en_mscbus;
wire      [4:0] DP0_31_in_mux_peripheral_mscbus;
wire      [1:0] DP0_31_out_demux_peripheral_mscbus;
wire            DP0_3_IO;
wire      [5:0] DP0_3_in_mux_en_mscbus;
wire      [5:0] DP0_3_in_mux_peripheral_mscbus;
wire      [1:0] DP0_3_out_demux_peripheral_mscbus;
wire            DP0_4_IO;
wire      [6:0] DP0_4_in_mux_en_mscbus;
wire      [6:0] DP0_4_in_mux_peripheral_mscbus;
wire            DP0_4_out_demux_peripheral_mscbus;
wire            DP0_5_IO;
wire      [5:0] DP0_5_in_mux_en_mscbus;
wire      [5:0] DP0_5_in_mux_peripheral_mscbus;
wire      [1:0] DP0_5_out_demux_peripheral_mscbus;
wire            DP0_6_IO;
wire      [6:0] DP0_6_in_mux_en_mscbus;
wire      [6:0] DP0_6_in_mux_peripheral_mscbus;
wire            DP0_6_out_demux_peripheral_mscbus;
wire            DP0_7_IO;
wire      [5:0] DP0_7_in_mux_en_mscbus;
wire      [5:0] DP0_7_in_mux_peripheral_mscbus;
wire      [1:0] DP0_7_out_demux_peripheral_mscbus;
wire            DP0_8_IO;
wire      [5:0] DP0_8_in_mux_en_mscbus;
wire      [5:0] DP0_8_in_mux_peripheral_mscbus;
wire      [1:0] DP0_8_out_demux_peripheral_mscbus;
wire            DP0_9_IO;
wire      [5:0] DP0_9_in_mux_en_mscbus;
wire      [5:0] DP0_9_in_mux_peripheral_mscbus;
wire      [1:0] DP0_9_out_demux_peripheral_mscbus;
wire            DP1_0_IO;
wire      [3:0] DP1_0_in_mux_en_mscbus;
wire      [3:0] DP1_0_in_mux_peripheral_mscbus;
wire      [2:0] DP1_0_out_demux_peripheral_mscbus;
wire            DP1_10_IO;
wire      [2:0] DP1_10_in_mux_en_mscbus;
wire      [2:0] DP1_10_in_mux_peripheral_mscbus;
wire      [2:0] DP1_10_out_demux_peripheral_mscbus;
wire            DP1_11_IO;
wire      [2:0] DP1_11_in_mux_en_mscbus;
wire      [2:0] DP1_11_in_mux_peripheral_mscbus;
wire      [2:0] DP1_11_out_demux_peripheral_mscbus;
wire            DP1_12_IO;
wire      [2:0] DP1_12_in_mux_en_mscbus;
wire      [2:0] DP1_12_in_mux_peripheral_mscbus;
wire      [1:0] DP1_12_out_demux_peripheral_mscbus;
wire            DP1_13_IO;
wire      [4:0] DP1_13_in_mux_en_mscbus;
wire      [4:0] DP1_13_in_mux_peripheral_mscbus;
wire      [1:0] DP1_13_out_demux_peripheral_mscbus;
wire            DP1_14_IO;
wire      [2:0] DP1_14_in_mux_en_mscbus;
wire      [2:0] DP1_14_in_mux_peripheral_mscbus;
wire      [3:0] DP1_14_out_demux_peripheral_mscbus;
wire            DP1_15_IO;
wire      [4:0] DP1_15_in_mux_en_mscbus;
wire      [4:0] DP1_15_in_mux_peripheral_mscbus;
wire      [1:0] DP1_15_out_demux_peripheral_mscbus;
wire            DP1_16_IO;
wire      [3:0] DP1_16_in_mux_en_mscbus;
wire      [3:0] DP1_16_in_mux_peripheral_mscbus;
wire      [2:0] DP1_16_out_demux_peripheral_mscbus;
wire            DP1_17_IO;
wire      [3:0] DP1_17_in_mux_en_mscbus;
wire      [3:0] DP1_17_in_mux_peripheral_mscbus;
wire      [2:0] DP1_17_out_demux_peripheral_mscbus;
wire            DP1_18_IO;
wire      [3:0] DP1_18_in_mux_en_mscbus;
wire      [3:0] DP1_18_in_mux_peripheral_mscbus;
wire      [2:0] DP1_18_out_demux_peripheral_mscbus;
wire            DP1_19_IO;
wire      [4:0] DP1_19_in_mux_en_mscbus;
wire      [4:0] DP1_19_in_mux_peripheral_mscbus;
wire      [1:0] DP1_19_out_demux_peripheral_mscbus;
wire            DP1_1_IO;
wire      [3:0] DP1_1_in_mux_en_mscbus;
wire      [3:0] DP1_1_in_mux_peripheral_mscbus;
wire      [2:0] DP1_1_out_demux_peripheral_mscbus;
wire            DP1_20_IO;
wire      [3:0] DP1_20_in_mux_en_mscbus;
wire      [3:0] DP1_20_in_mux_peripheral_mscbus;
wire      [2:0] DP1_20_out_demux_peripheral_mscbus;
wire            DP1_21_IO;
wire      [4:0] DP1_21_in_mux_en_mscbus;
wire      [4:0] DP1_21_in_mux_peripheral_mscbus;
wire      [1:0] DP1_21_out_demux_peripheral_mscbus;
wire            DP1_22_IO;
wire      [4:0] DP1_22_in_mux_en_mscbus;
wire      [4:0] DP1_22_in_mux_peripheral_mscbus;
wire      [1:0] DP1_22_out_demux_peripheral_mscbus;
wire            DP1_23_IO;
wire      [3:0] DP1_23_in_mux_en_mscbus;
wire      [3:0] DP1_23_in_mux_peripheral_mscbus;
wire      [1:0] DP1_23_out_demux_peripheral_mscbus;
wire            DP1_24_IO;
wire      [3:0] DP1_24_in_mux_en_mscbus;
wire      [3:0] DP1_24_in_mux_peripheral_mscbus;
wire      [1:0] DP1_24_out_demux_peripheral_mscbus;
wire            DP1_25_IO;
wire      [5:0] DP1_25_in_mux_en_mscbus;
wire      [5:0] DP1_25_in_mux_peripheral_mscbus;
wire            DP1_25_out_demux_peripheral_mscbus;
wire            DP1_26_IO;
wire      [5:0] DP1_26_in_mux_en_mscbus;
wire      [5:0] DP1_26_in_mux_peripheral_mscbus;
wire            DP1_26_out_demux_peripheral_mscbus;
wire            DP1_27_IO;
wire      [5:0] DP1_27_in_mux_en_mscbus;
wire      [5:0] DP1_27_in_mux_peripheral_mscbus;
wire            DP1_27_out_demux_peripheral_mscbus;
wire            DP1_28_IO;
wire      [4:0] DP1_28_in_mux_en_mscbus;
wire      [4:0] DP1_28_in_mux_peripheral_mscbus;
wire      [1:0] DP1_28_out_demux_peripheral_mscbus;
wire            DP1_29_IO;
wire      [4:0] DP1_29_in_mux_en_mscbus;
wire      [4:0] DP1_29_in_mux_peripheral_mscbus;
wire      [1:0] DP1_29_out_demux_peripheral_mscbus;
wire            DP1_2_IO;
wire      [3:0] DP1_2_in_mux_en_mscbus;
wire      [3:0] DP1_2_in_mux_peripheral_mscbus;
wire      [2:0] DP1_2_out_demux_peripheral_mscbus;
wire            DP1_30_IO;
wire      [4:0] DP1_30_in_mux_en_mscbus;
wire      [4:0] DP1_30_in_mux_peripheral_mscbus;
wire      [1:0] DP1_30_out_demux_peripheral_mscbus;
wire            DP1_31_IO;
wire      [3:0] DP1_31_in_mux_en_mscbus;
wire      [3:0] DP1_31_in_mux_peripheral_mscbus;
wire      [2:0] DP1_31_out_demux_peripheral_mscbus;
wire            DP1_3_IO;
wire      [4:0] DP1_3_in_mux_en_mscbus;
wire      [4:0] DP1_3_in_mux_peripheral_mscbus;
wire      [1:0] DP1_3_out_demux_peripheral_mscbus;
wire            DP1_4_IO;
wire      [4:0] DP1_4_in_mux_en_mscbus;
wire      [4:0] DP1_4_in_mux_peripheral_mscbus;
wire      [1:0] DP1_4_out_demux_peripheral_mscbus;
wire            DP1_5_IO;
wire      [4:0] DP1_5_in_mux_en_mscbus;
wire      [4:0] DP1_5_in_mux_peripheral_mscbus;
wire      [1:0] DP1_5_out_demux_peripheral_mscbus;
wire            DP1_6_IO;
wire      [3:0] DP1_6_in_mux_en_mscbus;
wire      [3:0] DP1_6_in_mux_peripheral_mscbus;
wire      [2:0] DP1_6_out_demux_peripheral_mscbus;
wire            DP1_7_IO;
wire      [4:0] DP1_7_in_mux_en_mscbus;
wire      [4:0] DP1_7_in_mux_peripheral_mscbus;
wire      [1:0] DP1_7_out_demux_peripheral_mscbus;
wire            DP1_8_IO;
wire      [3:0] DP1_8_in_mux_en_mscbus;
wire      [3:0] DP1_8_in_mux_peripheral_mscbus;
wire      [1:0] DP1_8_out_demux_peripheral_mscbus;
wire            DP1_9_IO;
wire      [3:0] DP1_9_in_mux_en_mscbus;
wire      [3:0] DP1_9_in_mux_peripheral_mscbus;
wire      [1:0] DP1_9_out_demux_peripheral_mscbus;
wire            DP2_0_IO;
wire      [4:0] DP2_0_in_mux_en_mscbus;
wire      [4:0] DP2_0_in_mux_peripheral_mscbus;
wire      [1:0] DP2_0_out_demux_peripheral_mscbus;
wire            DP2_10_IO;
wire      [4:0] DP2_10_in_mux_en_mscbus;
wire      [4:0] DP2_10_in_mux_peripheral_mscbus;
wire            DP2_10_out_demux_peripheral_mscbus;
wire            DP2_11_IO;
wire      [3:0] DP2_11_in_mux_en_mscbus;
wire      [3:0] DP2_11_in_mux_peripheral_mscbus;
wire            DP2_11_out_demux_peripheral_mscbus;
wire            DP2_12_IO;
wire      [4:0] DP2_12_in_mux_en_mscbus;
wire      [4:0] DP2_12_in_mux_peripheral_mscbus;
wire      [1:0] DP2_12_out_demux_peripheral_mscbus;
wire            DP2_13_IO;
wire      [5:0] DP2_13_in_mux_en_mscbus;
wire      [5:0] DP2_13_in_mux_peripheral_mscbus;
wire      [3:0] DP2_13_out_demux_peripheral_mscbus;
wire            DP2_14_IO;
wire      [6:0] DP2_14_in_mux_en_mscbus;
wire      [6:0] DP2_14_in_mux_peripheral_mscbus;
wire      [2:0] DP2_14_out_demux_peripheral_mscbus;
wire            DP2_15_IO;
wire      [5:0] DP2_15_in_mux_en_mscbus;
wire      [5:0] DP2_15_in_mux_peripheral_mscbus;
wire      [3:0] DP2_15_out_demux_peripheral_mscbus;
wire            DP2_16_IO;
wire      [5:0] DP2_16_in_mux_en_mscbus;
wire      [5:0] DP2_16_in_mux_peripheral_mscbus;
wire      [3:0] DP2_16_out_demux_peripheral_mscbus;
wire            DP2_17_IO;
wire      [5:0] DP2_17_in_mux_en_mscbus;
wire      [5:0] DP2_17_in_mux_peripheral_mscbus;
wire      [3:0] DP2_17_out_demux_peripheral_mscbus;
wire            DP2_18_IO;
wire      [6:0] DP2_18_in_mux_en_mscbus;
wire      [6:0] DP2_18_in_mux_peripheral_mscbus;
wire      [2:0] DP2_18_out_demux_peripheral_mscbus;
wire            DP2_19_IO;
wire      [6:0] DP2_19_in_mux_en_mscbus;
wire      [6:0] DP2_19_in_mux_peripheral_mscbus;
wire      [2:0] DP2_19_out_demux_peripheral_mscbus;
wire            DP2_1_IO;
wire      [4:0] DP2_1_in_mux_en_mscbus;
wire      [4:0] DP2_1_in_mux_peripheral_mscbus;
wire            DP2_1_out_demux_peripheral_mscbus;
wire            DP2_20_IO;
wire      [5:0] DP2_20_in_mux_en_mscbus;
wire      [5:0] DP2_20_in_mux_peripheral_mscbus;
wire      [3:0] DP2_20_out_demux_peripheral_mscbus;
wire            DP2_21_IO;
wire      [6:0] DP2_21_in_mux_en_mscbus;
wire      [6:0] DP2_21_in_mux_peripheral_mscbus;
wire            DP2_21_out_demux_peripheral_mscbus;
wire            DP2_22_IO;
wire      [5:0] DP2_22_in_mux_en_mscbus;
wire      [5:0] DP2_22_in_mux_peripheral_mscbus;
wire      [1:0] DP2_22_out_demux_peripheral_mscbus;
wire            DP2_23_IO;
wire      [6:0] DP2_23_in_mux_en_mscbus;
wire      [6:0] DP2_23_in_mux_peripheral_mscbus;
wire      [1:0] DP2_23_out_demux_peripheral_mscbus;
wire            DP2_24_IO;
wire      [5:0] DP2_24_in_mux_en_mscbus;
wire      [5:0] DP2_24_in_mux_peripheral_mscbus;
wire      [2:0] DP2_24_out_demux_peripheral_mscbus;
wire            DP2_25_IO;
wire      [6:0] DP2_25_in_mux_en_mscbus;
wire      [6:0] DP2_25_in_mux_peripheral_mscbus;
wire            DP2_25_out_demux_peripheral_mscbus;
wire            DP2_26_IO;
wire      [4:0] DP2_26_in_mux_en_mscbus;
wire      [4:0] DP2_26_in_mux_peripheral_mscbus;
wire      [2:0] DP2_26_out_demux_peripheral_mscbus;
wire            DP2_27_IO;
wire      [5:0] DP2_27_in_mux_en_mscbus;
wire      [5:0] DP2_27_in_mux_peripheral_mscbus;
wire      [1:0] DP2_27_out_demux_peripheral_mscbus;
wire            DP2_28_IO;
wire      [3:0] DP2_28_in_mux_en_mscbus;
wire      [3:0] DP2_28_in_mux_peripheral_mscbus;
wire      [3:0] DP2_28_out_demux_peripheral_mscbus;
wire            DP2_29_IO;
wire      [5:0] DP2_29_in_mux_en_mscbus;
wire      [5:0] DP2_29_in_mux_peripheral_mscbus;
wire      [1:0] DP2_29_out_demux_peripheral_mscbus;
wire            DP2_2_IO;
wire      [4:0] DP2_2_in_mux_en_mscbus;
wire      [4:0] DP2_2_in_mux_peripheral_mscbus;
wire      [1:0] DP2_2_out_demux_peripheral_mscbus;
wire            DP2_30_IO;
wire      [4:0] DP2_30_in_mux_en_mscbus;
wire      [4:0] DP2_30_in_mux_peripheral_mscbus;
wire      [2:0] DP2_30_out_demux_peripheral_mscbus;
wire            DP2_31_IO;
wire      [5:0] DP2_31_in_mux_en_mscbus;
wire      [5:0] DP2_31_in_mux_peripheral_mscbus;
wire      [1:0] DP2_31_out_demux_peripheral_mscbus;
wire            DP2_3_IO;
wire      [4:0] DP2_3_in_mux_en_mscbus;
wire      [4:0] DP2_3_in_mux_peripheral_mscbus;
wire      [1:0] DP2_3_out_demux_peripheral_mscbus;
wire            DP2_4_IO;
wire      [4:0] DP2_4_in_mux_en_mscbus;
wire      [4:0] DP2_4_in_mux_peripheral_mscbus;
wire            DP2_4_out_demux_peripheral_mscbus;
wire            DP2_5_IO;
wire      [4:0] DP2_5_in_mux_en_mscbus;
wire      [4:0] DP2_5_in_mux_peripheral_mscbus;
wire            DP2_5_out_demux_peripheral_mscbus;
wire            DP2_6_IO;
wire      [3:0] DP2_6_in_mux_en_mscbus;
wire      [3:0] DP2_6_in_mux_peripheral_mscbus;
wire      [1:0] DP2_6_out_demux_peripheral_mscbus;
wire            DP2_7_IO;
wire      [4:0] DP2_7_in_mux_en_mscbus;
wire      [4:0] DP2_7_in_mux_peripheral_mscbus;
wire            DP2_7_out_demux_peripheral_mscbus;
wire            DP2_8_IO;
wire      [4:0] DP2_8_in_mux_en_mscbus;
wire      [4:0] DP2_8_in_mux_peripheral_mscbus;
wire            DP2_8_out_demux_peripheral_mscbus;
wire            DP2_9_IO;
wire      [4:0] DP2_9_in_mux_en_mscbus;
wire      [4:0] DP2_9_in_mux_peripheral_mscbus;
wire            DP2_9_out_demux_peripheral_mscbus;
wire            DP3_0_IO;
wire      [4:0] DP3_0_in_mux_en_mscbus;
wire      [4:0] DP3_0_in_mux_peripheral_mscbus;
wire      [2:0] DP3_0_out_demux_peripheral_mscbus;
wire            DP3_10_IO;
wire      [3:0] DP3_10_in_mux_en_mscbus;
wire      [3:0] DP3_10_in_mux_peripheral_mscbus;
wire      [3:0] DP3_10_out_demux_peripheral_mscbus;
wire            DP3_11_IO;
wire      [4:0] DP3_11_in_mux_en_mscbus;
wire      [4:0] DP3_11_in_mux_peripheral_mscbus;
wire      [2:0] DP3_11_out_demux_peripheral_mscbus;
wire            DP3_12_IO;
wire      [6:0] DP3_12_in_mux_en_mscbus;
wire      [6:0] DP3_12_in_mux_peripheral_mscbus;
wire            DP3_12_out_demux_peripheral_mscbus;
wire            DP3_13_IO;
wire      [4:0] DP3_13_in_mux_en_mscbus;
wire      [4:0] DP3_13_in_mux_peripheral_mscbus;
wire      [2:0] DP3_13_out_demux_peripheral_mscbus;
wire            DP3_14_IO;
wire      [6:0] DP3_14_in_mux_en_mscbus;
wire      [6:0] DP3_14_in_mux_peripheral_mscbus;
wire            DP3_14_out_demux_peripheral_mscbus;
wire            DP3_15_IO;
wire      [5:0] DP3_15_in_mux_en_mscbus;
wire      [5:0] DP3_15_in_mux_peripheral_mscbus;
wire      [1:0] DP3_15_out_demux_peripheral_mscbus;
wire            DP3_16_IO;
wire      [5:0] DP3_16_in_mux_en_mscbus;
wire      [5:0] DP3_16_in_mux_peripheral_mscbus;
wire      [1:0] DP3_16_out_demux_peripheral_mscbus;
wire            DP3_17_IO;
wire      [4:0] DP3_17_in_mux_en_mscbus;
wire      [4:0] DP3_17_in_mux_peripheral_mscbus;
wire      [2:0] DP3_17_out_demux_peripheral_mscbus;
wire            DP3_18_IO;
wire      [6:0] DP3_18_in_mux_en_mscbus;
wire      [6:0] DP3_18_in_mux_peripheral_mscbus;
wire            DP3_18_out_demux_peripheral_mscbus;
wire            DP3_19_IO;
wire      [6:0] DP3_19_in_mux_en_mscbus;
wire      [6:0] DP3_19_in_mux_peripheral_mscbus;
wire            DP3_19_out_demux_peripheral_mscbus;
wire            DP3_1_IO;
wire      [4:0] DP3_1_in_mux_en_mscbus;
wire      [4:0] DP3_1_in_mux_peripheral_mscbus;
wire      [2:0] DP3_1_out_demux_peripheral_mscbus;
wire            DP3_20_IO;
wire      [6:0] DP3_20_in_mux_en_mscbus;
wire      [6:0] DP3_20_in_mux_peripheral_mscbus;
wire            DP3_20_out_demux_peripheral_mscbus;
wire            DP3_21_IO;
wire      [7:0] DP3_21_in_mux_en_mscbus;
wire      [7:0] DP3_21_in_mux_peripheral_mscbus;
wire            DP3_21_out_demux_peripheral_mscbus;
wire            DP3_22_IO;
wire      [7:0] DP3_22_in_mux_en_mscbus;
wire      [7:0] DP3_22_in_mux_peripheral_mscbus;
wire            DP3_22_out_demux_peripheral_mscbus;
wire            DP3_23_IO;
wire      [7:0] DP3_23_in_mux_en_mscbus;
wire      [7:0] DP3_23_in_mux_peripheral_mscbus;
wire            DP3_23_out_demux_peripheral_mscbus;
wire            DP3_24_IO;
wire      [5:0] DP3_24_in_mux_en_mscbus;
wire      [5:0] DP3_24_in_mux_peripheral_mscbus;
wire      [2:0] DP3_24_out_demux_peripheral_mscbus;
wire            DP3_25_IO;
wire      [6:0] DP3_25_in_mux_en_mscbus;
wire      [6:0] DP3_25_in_mux_peripheral_mscbus;
wire      [1:0] DP3_25_out_demux_peripheral_mscbus;
wire            DP3_26_IO;
wire      [5:0] DP3_26_in_mux_en_mscbus;
wire      [5:0] DP3_26_in_mux_peripheral_mscbus;
wire      [2:0] DP3_26_out_demux_peripheral_mscbus;
wire            DP3_27_IO;
wire      [4:0] DP3_27_in_mux_en_mscbus;
wire      [4:0] DP3_27_in_mux_peripheral_mscbus;
wire      [2:0] DP3_27_out_demux_peripheral_mscbus;
wire            DP3_28_IO;
wire      [5:0] DP3_28_in_mux_en_mscbus;
wire      [5:0] DP3_28_in_mux_peripheral_mscbus;
wire      [2:0] DP3_28_out_demux_peripheral_mscbus;
wire            DP3_29_IO;
wire      [6:0] DP3_29_in_mux_en_mscbus;
wire      [6:0] DP3_29_in_mux_peripheral_mscbus;
wire      [1:0] DP3_29_out_demux_peripheral_mscbus;
wire            DP3_2_IO;
wire      [5:0] DP3_2_in_mux_en_mscbus;
wire      [5:0] DP3_2_in_mux_peripheral_mscbus;
wire      [1:0] DP3_2_out_demux_peripheral_mscbus;
wire            DP3_30_IO;
wire      [6:0] DP3_30_in_mux_en_mscbus;
wire      [6:0] DP3_30_in_mux_peripheral_mscbus;
wire      [2:0] DP3_30_out_demux_peripheral_mscbus;
wire            DP3_31_IO;
wire      [4:0] DP3_31_in_mux_en_mscbus;
wire      [4:0] DP3_31_in_mux_peripheral_mscbus;
wire      [4:0] DP3_31_out_demux_peripheral_mscbus;
wire            DP3_3_IO;
wire      [3:0] DP3_3_in_mux_en_mscbus;
wire      [3:0] DP3_3_in_mux_peripheral_mscbus;
wire      [3:0] DP3_3_out_demux_peripheral_mscbus;
wire            DP3_4_IO;
wire      [5:0] DP3_4_in_mux_en_mscbus;
wire      [5:0] DP3_4_in_mux_peripheral_mscbus;
wire      [1:0] DP3_4_out_demux_peripheral_mscbus;
wire            DP3_5_IO;
wire      [4:0] DP3_5_in_mux_en_mscbus;
wire      [4:0] DP3_5_in_mux_peripheral_mscbus;
wire      [1:0] DP3_5_out_demux_peripheral_mscbus;
wire            DP3_6_IO;
wire      [4:0] DP3_6_in_mux_en_mscbus;
wire      [4:0] DP3_6_in_mux_peripheral_mscbus;
wire      [1:0] DP3_6_out_demux_peripheral_mscbus;
wire            DP3_7_IO;
wire      [4:0] DP3_7_in_mux_en_mscbus;
wire      [4:0] DP3_7_in_mux_peripheral_mscbus;
wire      [1:0] DP3_7_out_demux_peripheral_mscbus;
wire            DP3_8_IO;
wire      [5:0] DP3_8_in_mux_en_mscbus;
wire      [5:0] DP3_8_in_mux_peripheral_mscbus;
wire      [1:0] DP3_8_out_demux_peripheral_mscbus;
wire            DP3_9_IO;
wire      [4:0] DP3_9_in_mux_en_mscbus;
wire      [4:0] DP3_9_in_mux_peripheral_mscbus;
wire      [2:0] DP3_9_out_demux_peripheral_mscbus;
wire            DP4_0_IO;
wire      [5:0] DP4_0_in_mux_en_mscbus;
wire      [5:0] DP4_0_in_mux_peripheral_mscbus;
wire      [2:0] DP4_0_out_demux_peripheral_mscbus;
wire            DP4_10_IO;
wire      [6:0] DP4_10_in_mux_en_mscbus;
wire      [6:0] DP4_10_in_mux_peripheral_mscbus;
wire      [3:0] DP4_10_out_demux_peripheral_mscbus;
wire            DP4_11_IO;
wire      [7:0] DP4_11_in_mux_en_mscbus;
wire      [7:0] DP4_11_in_mux_peripheral_mscbus;
wire      [2:0] DP4_11_out_demux_peripheral_mscbus;
wire            DP4_12_IO;
wire      [6:0] DP4_12_in_mux_en_mscbus;
wire      [6:0] DP4_12_in_mux_peripheral_mscbus;
wire      [3:0] DP4_12_out_demux_peripheral_mscbus;
wire            DP4_13_IO;
wire      [6:0] DP4_13_in_mux_en_mscbus;
wire      [6:0] DP4_13_in_mux_peripheral_mscbus;
wire      [3:0] DP4_13_out_demux_peripheral_mscbus;
wire            DP4_14_IO;
wire      [5:0] DP4_14_in_mux_en_mscbus;
wire      [5:0] DP4_14_in_mux_peripheral_mscbus;
wire      [2:0] DP4_14_out_demux_peripheral_mscbus;
wire            DP4_15_IO;
wire      [4:0] DP4_15_in_mux_en_mscbus;
wire      [4:0] DP4_15_in_mux_peripheral_mscbus;
wire      [3:0] DP4_15_out_demux_peripheral_mscbus;
wire            DP4_16_IO;
wire      [4:0] DP4_16_in_mux_en_mscbus;
wire      [4:0] DP4_16_in_mux_peripheral_mscbus;
wire      [3:0] DP4_16_out_demux_peripheral_mscbus;
wire            DP4_17_IO;
wire      [4:0] DP4_17_in_mux_en_mscbus;
wire      [4:0] DP4_17_in_mux_peripheral_mscbus;
wire      [3:0] DP4_17_out_demux_peripheral_mscbus;
wire            DP4_18_IO;
wire      [2:0] DP4_18_in_mux_en_mscbus;
wire      [2:0] DP4_18_in_mux_peripheral_mscbus;
wire      [2:0] DP4_18_out_demux_peripheral_mscbus;
wire            DP4_19_IO;
wire      [4:0] DP4_19_in_mux_en_mscbus;
wire      [4:0] DP4_19_in_mux_peripheral_mscbus;
wire      [1:0] DP4_19_out_demux_peripheral_mscbus;
wire            DP4_1_IO;
wire      [4:0] DP4_1_in_mux_en_mscbus;
wire      [4:0] DP4_1_in_mux_peripheral_mscbus;
wire      [3:0] DP4_1_out_demux_peripheral_mscbus;
wire            DP4_20_IO;
wire      [7:0] DP4_20_in_mux_en_mscbus;
wire      [7:0] DP4_20_in_mux_peripheral_mscbus;
wire      [1:0] DP4_20_out_demux_peripheral_mscbus;
wire            DP4_21_IO;
wire      [7:0] DP4_21_in_mux_en_mscbus;
wire      [7:0] DP4_21_in_mux_peripheral_mscbus;
wire      [1:0] DP4_21_out_demux_peripheral_mscbus;
wire            DP4_22_IO;
wire      [6:0] DP4_22_in_mux_en_mscbus;
wire      [6:0] DP4_22_in_mux_peripheral_mscbus;
wire      [2:0] DP4_22_out_demux_peripheral_mscbus;
wire            DP4_23_IO;
wire      [7:0] DP4_23_in_mux_en_mscbus;
wire      [7:0] DP4_23_in_mux_peripheral_mscbus;
wire      [2:0] DP4_23_out_demux_peripheral_mscbus;
wire            DP4_24_IO;
wire      [7:0] DP4_24_in_mux_en_mscbus;
wire      [7:0] DP4_24_in_mux_peripheral_mscbus;
wire      [2:0] DP4_24_out_demux_peripheral_mscbus;
wire            DP4_25_IO;
wire      [5:0] DP4_25_in_mux_en_mscbus;
wire      [5:0] DP4_25_in_mux_peripheral_mscbus;
wire      [3:0] DP4_25_out_demux_peripheral_mscbus;
wire            DP4_26_IO;
wire      [6:0] DP4_26_in_mux_en_mscbus;
wire      [6:0] DP4_26_in_mux_peripheral_mscbus;
wire      [2:0] DP4_26_out_demux_peripheral_mscbus;
wire            DP4_27_IO;
wire      [5:0] DP4_27_in_mux_en_mscbus;
wire      [5:0] DP4_27_in_mux_peripheral_mscbus;
wire      [2:0] DP4_27_out_demux_peripheral_mscbus;
wire            DP4_28_IO;
wire      [6:0] DP4_28_in_mux_en_mscbus;
wire      [6:0] DP4_28_in_mux_peripheral_mscbus;
wire      [2:0] DP4_28_out_demux_peripheral_mscbus;
wire            DP4_29_IO;
wire      [5:0] DP4_29_in_mux_en_mscbus;
wire      [5:0] DP4_29_in_mux_peripheral_mscbus;
wire      [4:0] DP4_29_out_demux_peripheral_mscbus;
wire            DP4_2_IO;
wire      [5:0] DP4_2_in_mux_en_mscbus;
wire      [5:0] DP4_2_in_mux_peripheral_mscbus;
wire      [2:0] DP4_2_out_demux_peripheral_mscbus;
wire            DP4_30_IO;
wire      [5:0] DP4_30_in_mux_en_mscbus;
wire      [5:0] DP4_30_in_mux_peripheral_mscbus;
wire      [2:0] DP4_30_out_demux_peripheral_mscbus;
wire            DP4_31_IO;
wire      [4:0] DP4_31_in_mux_en_mscbus;
wire      [4:0] DP4_31_in_mux_peripheral_mscbus;
wire      [3:0] DP4_31_out_demux_peripheral_mscbus;
wire            DP4_3_IO;
wire      [5:0] DP4_3_in_mux_en_mscbus;
wire      [5:0] DP4_3_in_mux_peripheral_mscbus;
wire      [2:0] DP4_3_out_demux_peripheral_mscbus;
wire            DP4_4_IO;
wire      [4:0] DP4_4_in_mux_en_mscbus;
wire      [4:0] DP4_4_in_mux_peripheral_mscbus;
wire      [3:0] DP4_4_out_demux_peripheral_mscbus;
wire            DP4_5_IO;
wire      [5:0] DP4_5_in_mux_en_mscbus;
wire      [5:0] DP4_5_in_mux_peripheral_mscbus;
wire            DP4_5_out_demux_peripheral_mscbus;
wire            DP4_6_IO;
wire      [6:0] DP4_6_in_mux_en_mscbus;
wire      [6:0] DP4_6_in_mux_peripheral_mscbus;
wire      [2:0] DP4_6_out_demux_peripheral_mscbus;
wire            DP4_7_IO;
wire      [7:0] DP4_7_in_mux_en_mscbus;
wire      [7:0] DP4_7_in_mux_peripheral_mscbus;
wire      [2:0] DP4_7_out_demux_peripheral_mscbus;
wire            DP4_8_IO;
wire      [8:0] DP4_8_in_mux_en_mscbus;
wire      [8:0] DP4_8_in_mux_peripheral_mscbus;
wire      [1:0] DP4_8_out_demux_peripheral_mscbus;
wire            DP4_9_IO;
wire      [6:0] DP4_9_in_mux_en_mscbus;
wire      [6:0] DP4_9_in_mux_peripheral_mscbus;
wire      [3:0] DP4_9_out_demux_peripheral_mscbus;
wire            DP5_0_IO;
wire      [7:0] DP5_0_in_mux_en_mscbus;
wire      [7:0] DP5_0_in_mux_peripheral_mscbus;
wire            DP5_0_out_demux_peripheral_mscbus;
wire            DP5_10_IO;
wire      [5:0] DP5_10_in_mux_en_mscbus;
wire      [5:0] DP5_10_in_mux_peripheral_mscbus;
wire      [2:0] DP5_10_out_demux_peripheral_mscbus;
wire            DP5_11_IO;
wire      [4:0] DP5_11_in_mux_en_mscbus;
wire      [4:0] DP5_11_in_mux_peripheral_mscbus;
wire      [3:0] DP5_11_out_demux_peripheral_mscbus;
wire            DP5_12_IO;
wire      [5:0] DP5_12_in_mux_en_mscbus;
wire      [5:0] DP5_12_in_mux_peripheral_mscbus;
wire      [2:0] DP5_12_out_demux_peripheral_mscbus;
wire            DP5_13_IO;
wire      [5:0] DP5_13_in_mux_en_mscbus;
wire      [5:0] DP5_13_in_mux_peripheral_mscbus;
wire      [2:0] DP5_13_out_demux_peripheral_mscbus;
wire            DP5_14_IO;
wire      [6:0] DP5_14_in_mux_en_mscbus;
wire      [6:0] DP5_14_in_mux_peripheral_mscbus;
wire            DP5_14_out_demux_peripheral_mscbus;
wire            DP5_15_IO;
wire      [5:0] DP5_15_in_mux_en_mscbus;
wire      [5:0] DP5_15_in_mux_peripheral_mscbus;
wire      [1:0] DP5_15_out_demux_peripheral_mscbus;
wire            DP5_16_IO;
wire      [5:0] DP5_16_in_mux_en_mscbus;
wire      [5:0] DP5_16_in_mux_peripheral_mscbus;
wire      [1:0] DP5_16_out_demux_peripheral_mscbus;
wire            DP5_17_IO;
wire      [5:0] DP5_17_in_mux_en_mscbus;
wire      [5:0] DP5_17_in_mux_peripheral_mscbus;
wire      [1:0] DP5_17_out_demux_peripheral_mscbus;
wire            DP5_18_IO;
wire      [5:0] DP5_18_in_mux_en_mscbus;
wire      [5:0] DP5_18_in_mux_peripheral_mscbus;
wire            DP5_18_out_demux_peripheral_mscbus;
wire            DP5_19_IO;
wire      [4:0] DP5_19_in_mux_en_mscbus;
wire      [4:0] DP5_19_in_mux_peripheral_mscbus;
wire      [1:0] DP5_19_out_demux_peripheral_mscbus;
wire            DP5_1_IO;
wire      [6:0] DP5_1_in_mux_en_mscbus;
wire      [6:0] DP5_1_in_mux_peripheral_mscbus;
wire      [2:0] DP5_1_out_demux_peripheral_mscbus;
wire            DP5_20_IO;
wire      [6:0] DP5_20_in_mux_en_mscbus;
wire      [6:0] DP5_20_in_mux_peripheral_mscbus;
wire            DP5_20_out_demux_peripheral_mscbus;
wire            DP5_21_IO;
wire      [5:0] DP5_21_in_mux_en_mscbus;
wire      [5:0] DP5_21_in_mux_peripheral_mscbus;
wire      [1:0] DP5_21_out_demux_peripheral_mscbus;
wire            DP5_22_IO;
wire      [4:0] DP5_22_in_mux_en_mscbus;
wire      [4:0] DP5_22_in_mux_peripheral_mscbus;
wire      [2:0] DP5_22_out_demux_peripheral_mscbus;
wire            DP5_23_IO;
wire      [5:0] DP5_23_in_mux_en_mscbus;
wire      [5:0] DP5_23_in_mux_peripheral_mscbus;
wire      [1:0] DP5_23_out_demux_peripheral_mscbus;
wire            DP5_24_IO;
wire      [5:0] DP5_24_in_mux_en_mscbus;
wire      [5:0] DP5_24_in_mux_peripheral_mscbus;
wire      [1:0] DP5_24_out_demux_peripheral_mscbus;
wire            DP5_25_IO;
wire      [4:0] DP5_25_in_mux_en_mscbus;
wire      [4:0] DP5_25_in_mux_peripheral_mscbus;
wire      [1:0] DP5_25_out_demux_peripheral_mscbus;
wire            DP5_26_IO;
wire      [6:0] DP5_26_in_mux_en_mscbus;
wire      [6:0] DP5_26_in_mux_peripheral_mscbus;
wire      [1:0] DP5_26_out_demux_peripheral_mscbus;
wire            DP5_27_IO;
wire      [8:0] DP5_27_in_mux_en_mscbus;
wire      [8:0] DP5_27_in_mux_peripheral_mscbus;
wire            DP5_27_out_demux_peripheral_mscbus;
wire            DP5_28_IO;
wire      [6:0] DP5_28_in_mux_en_mscbus;
wire      [6:0] DP5_28_in_mux_peripheral_mscbus;
wire      [2:0] DP5_28_out_demux_peripheral_mscbus;
wire            DP5_29_IO;
wire      [7:0] DP5_29_in_mux_en_mscbus;
wire      [7:0] DP5_29_in_mux_peripheral_mscbus;
wire      [1:0] DP5_29_out_demux_peripheral_mscbus;
wire            DP5_2_IO;
wire      [5:0] DP5_2_in_mux_en_mscbus;
wire      [5:0] DP5_2_in_mux_peripheral_mscbus;
wire      [1:0] DP5_2_out_demux_peripheral_mscbus;
wire            DP5_30_IO;
wire      [5:0] DP5_30_in_mux_en_mscbus;
wire      [5:0] DP5_30_in_mux_peripheral_mscbus;
wire      [3:0] DP5_30_out_demux_peripheral_mscbus;
wire            DP5_31_IO;
wire      [7:0] DP5_31_in_mux_en_mscbus;
wire      [7:0] DP5_31_in_mux_peripheral_mscbus;
wire      [1:0] DP5_31_out_demux_peripheral_mscbus;
wire            DP5_3_IO;
wire      [5:0] DP5_3_in_mux_en_mscbus;
wire      [5:0] DP5_3_in_mux_peripheral_mscbus;
wire      [1:0] DP5_3_out_demux_peripheral_mscbus;
wire            DP5_4_IO;
wire      [5:0] DP5_4_in_mux_en_mscbus;
wire      [5:0] DP5_4_in_mux_peripheral_mscbus;
wire      [2:0] DP5_4_out_demux_peripheral_mscbus;
wire            DP5_5_IO;
wire      [5:0] DP5_5_in_mux_en_mscbus;
wire      [5:0] DP5_5_in_mux_peripheral_mscbus;
wire      [2:0] DP5_5_out_demux_peripheral_mscbus;
wire            DP5_6_IO;
wire      [7:0] DP5_6_in_mux_en_mscbus;
wire      [7:0] DP5_6_in_mux_peripheral_mscbus;
wire      [1:0] DP5_6_out_demux_peripheral_mscbus;
wire            DP5_7_IO;
wire      [7:0] DP5_7_in_mux_en_mscbus;
wire      [7:0] DP5_7_in_mux_peripheral_mscbus;
wire            DP5_7_out_demux_peripheral_mscbus;
wire            DP5_8_IO;
wire      [6:0] DP5_8_in_mux_en_mscbus;
wire      [6:0] DP5_8_in_mux_peripheral_mscbus;
wire      [1:0] DP5_8_out_demux_peripheral_mscbus;
wire            DP5_9_IO;
wire      [3:0] DP5_9_in_mux_en_mscbus;
wire      [3:0] DP5_9_in_mux_peripheral_mscbus;
wire      [4:0] DP5_9_out_demux_peripheral_mscbus;
wire            DP6_0_IO;
wire      [5:0] DP6_0_in_mux_en_mscbus;
wire      [5:0] DP6_0_in_mux_peripheral_mscbus;
wire      [3:0] DP6_0_out_demux_peripheral_mscbus;
wire            DP6_10_IO;
wire      [6:0] DP6_10_in_mux_en_mscbus;
wire      [6:0] DP6_10_in_mux_peripheral_mscbus;
wire      [2:0] DP6_10_out_demux_peripheral_mscbus;
wire            DP6_11_IO;
wire      [7:0] DP6_11_in_mux_en_mscbus;
wire      [7:0] DP6_11_in_mux_peripheral_mscbus;
wire      [1:0] DP6_11_out_demux_peripheral_mscbus;
wire            DP6_12_IO;
wire      [6:0] DP6_12_in_mux_en_mscbus;
wire      [6:0] DP6_12_in_mux_peripheral_mscbus;
wire      [1:0] DP6_12_out_demux_peripheral_mscbus;
wire            DP6_13_IO;
wire      [6:0] DP6_13_in_mux_en_mscbus;
wire      [6:0] DP6_13_in_mux_peripheral_mscbus;
wire      [2:0] DP6_13_out_demux_peripheral_mscbus;
wire            DP6_14_IO;
wire      [6:0] DP6_14_in_mux_en_mscbus;
wire      [6:0] DP6_14_in_mux_peripheral_mscbus;
wire      [1:0] DP6_14_out_demux_peripheral_mscbus;
wire            DP6_15_IO;
wire      [5:0] DP6_15_in_mux_en_mscbus;
wire      [5:0] DP6_15_in_mux_peripheral_mscbus;
wire      [2:0] DP6_15_out_demux_peripheral_mscbus;
wire            DP6_16_IO;
wire      [6:0] DP6_16_in_mux_en_mscbus;
wire      [6:0] DP6_16_in_mux_peripheral_mscbus;
wire      [1:0] DP6_16_out_demux_peripheral_mscbus;
wire            DP6_17_IO;
wire      [7:0] DP6_17_in_mux_en_mscbus;
wire      [7:0] DP6_17_in_mux_peripheral_mscbus;
wire            DP6_17_out_demux_peripheral_mscbus;
wire            DP6_18_IO;
wire      [7:0] DP6_18_in_mux_en_mscbus;
wire      [7:0] DP6_18_in_mux_peripheral_mscbus;
wire      [1:0] DP6_18_out_demux_peripheral_mscbus;
wire            DP6_19_IO;
wire      [5:0] DP6_19_in_mux_en_mscbus;
wire      [5:0] DP6_19_in_mux_peripheral_mscbus;
wire      [2:0] DP6_19_out_demux_peripheral_mscbus;
wire            DP6_1_IO;
wire      [5:0] DP6_1_in_mux_en_mscbus;
wire      [5:0] DP6_1_in_mux_peripheral_mscbus;
wire      [2:0] DP6_1_out_demux_peripheral_mscbus;
wire            DP6_20_IO;
wire      [7:0] DP6_20_in_mux_en_mscbus;
wire      [7:0] DP6_20_in_mux_peripheral_mscbus;
wire            DP6_20_out_demux_peripheral_mscbus;
wire            DP6_21_IO;
wire      [4:0] DP6_21_in_mux_en_mscbus;
wire      [4:0] DP6_21_in_mux_peripheral_mscbus;
wire      [3:0] DP6_21_out_demux_peripheral_mscbus;
wire            DP6_22_IO;
wire      [5:0] DP6_22_in_mux_en_mscbus;
wire      [5:0] DP6_22_in_mux_peripheral_mscbus;
wire      [2:0] DP6_22_out_demux_peripheral_mscbus;
wire            DP6_23_IO;
wire      [6:0] DP6_23_in_mux_en_mscbus;
wire      [6:0] DP6_23_in_mux_peripheral_mscbus;
wire      [1:0] DP6_23_out_demux_peripheral_mscbus;
wire            DP6_24_IO;
wire      [6:0] DP6_24_in_mux_en_mscbus;
wire      [6:0] DP6_24_in_mux_peripheral_mscbus;
wire      [1:0] DP6_24_out_demux_peripheral_mscbus;
wire            DP6_25_IO;
wire      [5:0] DP6_25_in_mux_en_mscbus;
wire      [5:0] DP6_25_in_mux_peripheral_mscbus;
wire      [2:0] DP6_25_out_demux_peripheral_mscbus;
wire            DP6_26_IO;
wire      [5:0] DP6_26_in_mux_en_mscbus;
wire      [5:0] DP6_26_in_mux_peripheral_mscbus;
wire            DP6_26_out_demux_peripheral_mscbus;
wire            DP6_27_IO;
wire      [5:0] DP6_27_in_mux_en_mscbus;
wire      [5:0] DP6_27_in_mux_peripheral_mscbus;
wire      [2:0] DP6_27_out_demux_peripheral_mscbus;
wire            DP6_2_IO;
wire      [5:0] DP6_2_in_mux_en_mscbus;
wire      [5:0] DP6_2_in_mux_peripheral_mscbus;
wire      [3:0] DP6_2_out_demux_peripheral_mscbus;
wire            DP6_3_IO;
wire      [7:0] DP6_3_in_mux_en_mscbus;
wire      [7:0] DP6_3_in_mux_peripheral_mscbus;
wire      [1:0] DP6_3_out_demux_peripheral_mscbus;
wire            DP6_4_IO;
wire      [5:0] DP6_4_in_mux_en_mscbus;
wire      [5:0] DP6_4_in_mux_peripheral_mscbus;
wire      [2:0] DP6_4_out_demux_peripheral_mscbus;
wire            DP6_5_IO;
wire      [5:0] DP6_5_in_mux_en_mscbus;
wire      [5:0] DP6_5_in_mux_peripheral_mscbus;
wire      [2:0] DP6_5_out_demux_peripheral_mscbus;
wire            DP6_6_IO;
wire      [7:0] DP6_6_in_mux_en_mscbus;
wire      [7:0] DP6_6_in_mux_peripheral_mscbus;
wire      [2:0] DP6_6_out_demux_peripheral_mscbus;
wire            DP6_7_IO;
wire      [7:0] DP6_7_in_mux_en_mscbus;
wire      [7:0] DP6_7_in_mux_peripheral_mscbus;
wire      [2:0] DP6_7_out_demux_peripheral_mscbus;
wire            DP6_8_IO;
wire      [5:0] DP6_8_in_mux_en_mscbus;
wire      [5:0] DP6_8_in_mux_peripheral_mscbus;
wire      [3:0] DP6_8_out_demux_peripheral_mscbus;
wire            DP6_9_IO;
wire      [6:0] DP6_9_in_mux_en_mscbus;
wire      [6:0] DP6_9_in_mux_peripheral_mscbus;
wire      [2:0] DP6_9_out_demux_peripheral_mscbus;
wire            DP7_0_IO;
wire      [6:0] DP7_0_in_mux_en_mscbus;
wire      [6:0] DP7_0_in_mux_peripheral_mscbus;
wire            DP7_0_out_demux_peripheral_mscbus;
wire            DP7_10_IO;
wire      [1:0] DP7_10_in_mux_en_mscbus;
wire      [1:0] DP7_10_in_mux_peripheral_mscbus;
wire      [3:0] DP7_10_out_demux_peripheral_mscbus;
wire            DP7_11_IO;
wire      [3:0] DP7_11_in_mux_en_mscbus;
wire      [3:0] DP7_11_in_mux_peripheral_mscbus;
wire      [1:0] DP7_11_out_demux_peripheral_mscbus;
wire            DP7_12_IO;
wire      [2:0] DP7_12_in_mux_en_mscbus;
wire      [2:0] DP7_12_in_mux_peripheral_mscbus;
wire      [2:0] DP7_12_out_demux_peripheral_mscbus;
wire            DP7_13_IO;
wire      [2:0] DP7_13_in_mux_en_mscbus;
wire      [2:0] DP7_13_in_mux_peripheral_mscbus;
wire      [2:0] DP7_13_out_demux_peripheral_mscbus;
wire            DP7_14_IO;
wire      [1:0] DP7_14_in_mux_en_mscbus;
wire      [1:0] DP7_14_in_mux_peripheral_mscbus;
wire      [3:0] DP7_14_out_demux_peripheral_mscbus;
wire            DP7_15_IO;
wire      [1:0] DP7_15_in_mux_en_mscbus;
wire      [1:0] DP7_15_in_mux_peripheral_mscbus;
wire      [2:0] DP7_15_out_demux_peripheral_mscbus;
wire            DP7_1_IO;
wire      [4:0] DP7_1_in_mux_en_mscbus;
wire      [4:0] DP7_1_in_mux_peripheral_mscbus;
wire      [2:0] DP7_1_out_demux_peripheral_mscbus;
wire            DP7_2_IO;
wire      [6:0] DP7_2_in_mux_en_mscbus;
wire      [6:0] DP7_2_in_mux_peripheral_mscbus;
wire            DP7_2_out_demux_peripheral_mscbus;
wire            DP7_3_IO;
wire      [6:0] DP7_3_in_mux_en_mscbus;
wire      [6:0] DP7_3_in_mux_peripheral_mscbus;
wire            DP7_3_out_demux_peripheral_mscbus;
wire            DP7_4_IO;
wire      [6:0] DP7_4_in_mux_en_mscbus;
wire      [6:0] DP7_4_in_mux_peripheral_mscbus;
wire            DP7_4_out_demux_peripheral_mscbus;
wire            DP7_5_IO;
wire      [6:0] DP7_5_in_mux_en_mscbus;
wire      [6:0] DP7_5_in_mux_peripheral_mscbus;
wire            DP7_5_out_demux_peripheral_mscbus;
wire            DP7_6_IO;
wire      [5:0] DP7_6_in_mux_en_mscbus;
wire      [5:0] DP7_6_in_mux_peripheral_mscbus;
wire      [1:0] DP7_6_out_demux_peripheral_mscbus;
wire            DP7_7_IO;
wire      [5:0] DP7_7_in_mux_en_mscbus;
wire      [5:0] DP7_7_in_mux_peripheral_mscbus;
wire      [2:0] DP7_7_out_demux_peripheral_mscbus;
wire            DP7_8_IO;
wire      [6:0] DP7_8_in_mux_en_mscbus;
wire      [6:0] DP7_8_in_mux_peripheral_mscbus;
wire      [1:0] DP7_8_out_demux_peripheral_mscbus;
wire            DP7_9_IO;
wire      [6:0] DP7_9_in_mux_en_mscbus;
wire      [6:0] DP7_9_in_mux_peripheral_mscbus;
wire      [2:0] DP7_9_out_demux_peripheral_mscbus;
wire            ERROR_IO;
wire            EXTPMICEN_IO;
wire            FLASHTESTPAD1FT_IO;
wire            FLASHTESTPAD2_IO;
wire            FLASHTESTPAD3FT_IO;
wire            FLASHTESTPAD4_IO;
wire            FLASHTESTPAD5_IO;
wire            MP0_0_IO;
wire      [3:0] MP0_0_in_mux_en_mscbus;
wire      [3:0] MP0_0_in_mux_peripheral_mscbus;
wire      [1:0] MP0_0_out_demux_peripheral_mscbus;
wire            MP0_10_IO;
wire      [3:0] MP0_10_in_mux_en_mscbus;
wire      [3:0] MP0_10_in_mux_peripheral_mscbus;
wire      [1:0] MP0_10_out_demux_peripheral_mscbus;
wire            MP0_11_IO;
wire            MP0_11_in_mux_en_mscbus;
wire            MP0_11_in_mux_peripheral_mscbus;
wire      [3:0] MP0_11_out_demux_peripheral_mscbus;
wire            MP0_12_IO;
wire      [3:0] MP0_12_in_mux_en_mscbus;
wire      [3:0] MP0_12_in_mux_peripheral_mscbus;
wire      [1:0] MP0_12_out_demux_peripheral_mscbus;
wire            MP0_13_IO;
wire      [1:0] MP0_13_in_mux_en_mscbus;
wire      [1:0] MP0_13_in_mux_peripheral_mscbus;
wire      [3:0] MP0_13_out_demux_peripheral_mscbus;
wire            MP0_14_IO;
wire      [4:0] MP0_14_in_mux_en_mscbus;
wire      [4:0] MP0_14_in_mux_peripheral_mscbus;
wire            MP0_14_out_demux_peripheral_mscbus;
wire            MP0_15_IO;
wire      [2:0] MP0_15_in_mux_en_mscbus;
wire      [2:0] MP0_15_in_mux_peripheral_mscbus;
wire      [2:0] MP0_15_out_demux_peripheral_mscbus;
wire            MP0_16_IO;
wire      [4:0] MP0_16_in_mux_en_mscbus;
wire      [4:0] MP0_16_in_mux_peripheral_mscbus;
wire            MP0_16_out_demux_peripheral_mscbus;
wire            MP0_17_IO;
wire            MP0_17_in_mux_en_mscbus;
wire            MP0_17_in_mux_peripheral_mscbus;
wire      [2:0] MP0_17_out_demux_peripheral_mscbus;
wire            MP0_18_IO;
wire      [4:0] MP0_18_in_mux_en_mscbus;
wire      [4:0] MP0_18_in_mux_peripheral_mscbus;
wire            MP0_18_out_demux_peripheral_mscbus;
wire            MP0_19_IO;
wire      [2:0] MP0_19_in_mux_en_mscbus;
wire      [2:0] MP0_19_in_mux_peripheral_mscbus;
wire      [2:0] MP0_19_out_demux_peripheral_mscbus;
wire            MP0_1_IO;
wire      [2:0] MP0_1_in_mux_en_mscbus;
wire      [2:0] MP0_1_in_mux_peripheral_mscbus;
wire      [2:0] MP0_1_out_demux_peripheral_mscbus;
wire            MP0_20_IO;
wire      [4:0] MP0_20_in_mux_en_mscbus;
wire      [4:0] MP0_20_in_mux_peripheral_mscbus;
wire            MP0_20_out_demux_peripheral_mscbus;
wire            MP0_21_IO;
wire      [2:0] MP0_21_in_mux_en_mscbus;
wire      [2:0] MP0_21_in_mux_peripheral_mscbus;
wire      [2:0] MP0_21_out_demux_peripheral_mscbus;
wire            MP0_22_IO;
wire      [3:0] MP0_22_in_mux_en_mscbus;
wire      [3:0] MP0_22_in_mux_peripheral_mscbus;
wire            MP0_22_out_demux_peripheral_mscbus;
wire            MP0_23_IO;
wire      [1:0] MP0_23_in_mux_en_mscbus;
wire      [1:0] MP0_23_in_mux_peripheral_mscbus;
wire      [1:0] MP0_23_out_demux_peripheral_mscbus;
wire            MP0_24_IO;
wire      [2:0] MP0_24_in_mux_en_mscbus;
wire      [2:0] MP0_24_in_mux_peripheral_mscbus;
wire      [3:0] MP0_24_out_demux_peripheral_mscbus;
wire            MP0_25_IO;
wire      [1:0] MP0_25_in_mux_en_mscbus;
wire      [1:0] MP0_25_in_mux_peripheral_mscbus;
wire      [4:0] MP0_25_out_demux_peripheral_mscbus;
wire            MP0_26_IO;
wire      [3:0] MP0_26_in_mux_en_mscbus;
wire      [3:0] MP0_26_in_mux_peripheral_mscbus;
wire      [2:0] MP0_26_out_demux_peripheral_mscbus;
wire            MP0_27_IO;
wire      [1:0] MP0_27_in_mux_en_mscbus;
wire      [1:0] MP0_27_in_mux_peripheral_mscbus;
wire      [4:0] MP0_27_out_demux_peripheral_mscbus;
wire            MP0_28_IO;
wire      [3:0] MP0_28_in_mux_en_mscbus;
wire      [3:0] MP0_28_in_mux_peripheral_mscbus;
wire            MP0_28_out_demux_peripheral_mscbus;
wire            MP0_29_IO;
wire            MP0_29_in_mux_en_mscbus;
wire            MP0_29_in_mux_peripheral_mscbus;
wire      [2:0] MP0_29_out_demux_peripheral_mscbus;
wire            MP0_2_IO;
wire      [3:0] MP0_2_in_mux_en_mscbus;
wire      [3:0] MP0_2_in_mux_peripheral_mscbus;
wire      [1:0] MP0_2_out_demux_peripheral_mscbus;
wire            MP0_30_IO;
wire      [4:0] MP0_30_in_mux_en_mscbus;
wire      [4:0] MP0_30_in_mux_peripheral_mscbus;
wire      [1:0] MP0_30_out_demux_peripheral_mscbus;
wire            MP0_31_IO;
wire      [3:0] MP0_31_in_mux_en_mscbus;
wire      [3:0] MP0_31_in_mux_peripheral_mscbus;
wire      [2:0] MP0_31_out_demux_peripheral_mscbus;
wire            MP0_3_IO;
wire      [2:0] MP0_3_in_mux_en_mscbus;
wire      [2:0] MP0_3_in_mux_peripheral_mscbus;
wire      [2:0] MP0_3_out_demux_peripheral_mscbus;
wire            MP0_4_IO;
wire      [3:0] MP0_4_in_mux_en_mscbus;
wire      [3:0] MP0_4_in_mux_peripheral_mscbus;
wire      [1:0] MP0_4_out_demux_peripheral_mscbus;
wire            MP0_5_IO;
wire            MP0_5_in_mux_en_mscbus;
wire            MP0_5_in_mux_peripheral_mscbus;
wire      [2:0] MP0_5_out_demux_peripheral_mscbus;
wire            MP0_6_IO;
wire      [3:0] MP0_6_in_mux_en_mscbus;
wire      [3:0] MP0_6_in_mux_peripheral_mscbus;
wire      [1:0] MP0_6_out_demux_peripheral_mscbus;
wire            MP0_7_IO;
wire      [2:0] MP0_7_in_mux_en_mscbus;
wire      [2:0] MP0_7_in_mux_peripheral_mscbus;
wire      [2:0] MP0_7_out_demux_peripheral_mscbus;
wire            MP0_8_IO;
wire      [4:0] MP0_8_in_mux_en_mscbus;
wire      [4:0] MP0_8_in_mux_peripheral_mscbus;
wire      [1:0] MP0_8_out_demux_peripheral_mscbus;
wire            MP0_9_IO;
wire      [1:0] MP0_9_in_mux_en_mscbus;
wire      [1:0] MP0_9_in_mux_peripheral_mscbus;
wire      [3:0] MP0_9_out_demux_peripheral_mscbus;
wire            MP1_0_IO;
wire      [4:0] MP1_0_in_mux_en_mscbus;
wire      [4:0] MP1_0_in_mux_peripheral_mscbus;
wire      [1:0] MP1_0_out_demux_peripheral_mscbus;
wire            MP1_10_IO;
wire      [2:0] MP1_10_in_mux_en_mscbus;
wire      [2:0] MP1_10_in_mux_peripheral_mscbus;
wire            MP1_10_out_demux_peripheral_mscbus;
wire            MP1_11_IO;
wire      [2:0] MP1_11_in_mux_en_mscbus;
wire      [2:0] MP1_11_in_mux_peripheral_mscbus;
wire            MP1_11_out_demux_peripheral_mscbus;
wire            MP1_12_IO;
wire      [1:0] MP1_12_in_mux_en_mscbus;
wire      [1:0] MP1_12_in_mux_peripheral_mscbus;
wire            MP1_12_out_demux_peripheral_mscbus;
wire            MP1_13_IO;
wire      [1:0] MP1_13_in_mux_en_mscbus;
wire      [1:0] MP1_13_in_mux_peripheral_mscbus;
wire            MP1_13_out_demux_peripheral_mscbus;
wire            MP1_14_IO;
wire      [1:0] MP1_14_in_mux_en_mscbus;
wire      [1:0] MP1_14_in_mux_peripheral_mscbus;
wire            MP1_14_out_demux_peripheral_mscbus;
wire            MP1_15_IO;
wire      [1:0] MP1_15_in_mux_en_mscbus;
wire      [1:0] MP1_15_in_mux_peripheral_mscbus;
wire            MP1_15_out_demux_peripheral_mscbus;
wire            MP1_1_IO;
wire      [3:0] MP1_1_in_mux_en_mscbus;
wire      [3:0] MP1_1_in_mux_peripheral_mscbus;
wire      [2:0] MP1_1_out_demux_peripheral_mscbus;
wire            MP1_2_IO;
wire      [2:0] MP1_2_in_mux_en_mscbus;
wire      [2:0] MP1_2_in_mux_peripheral_mscbus;
wire      [1:0] MP1_2_out_demux_peripheral_mscbus;
wire            MP1_3_IO;
wire            MP1_3_in_mux_en_mscbus;
wire            MP1_3_in_mux_peripheral_mscbus;
wire      [2:0] MP1_3_out_demux_peripheral_mscbus;
wire            MP1_4_IO;
wire      [1:0] MP1_4_in_mux_en_mscbus;
wire      [1:0] MP1_4_in_mux_peripheral_mscbus;
wire      [1:0] MP1_4_out_demux_peripheral_mscbus;
wire            MP1_5_IO;
wire      [1:0] MP1_5_in_mux_en_mscbus;
wire      [1:0] MP1_5_in_mux_peripheral_mscbus;
wire      [1:0] MP1_5_out_demux_peripheral_mscbus;
wire            MP1_6_IO;
wire      [1:0] MP1_6_in_mux_en_mscbus;
wire      [1:0] MP1_6_in_mux_peripheral_mscbus;
wire      [1:0] MP1_6_out_demux_peripheral_mscbus;
wire            MP1_7_IO;
wire      [1:0] MP1_7_in_mux_en_mscbus;
wire      [1:0] MP1_7_in_mux_peripheral_mscbus;
wire      [1:0] MP1_7_out_demux_peripheral_mscbus;
wire            MP1_8_IO;
wire      [1:0] MP1_8_in_mux_en_mscbus;
wire      [1:0] MP1_8_in_mux_peripheral_mscbus;
wire      [1:0] MP1_8_out_demux_peripheral_mscbus;
wire            MP1_9_IO;
wire      [1:0] MP1_9_in_mux_en_mscbus;
wire      [1:0] MP1_9_in_mux_peripheral_mscbus;
wire      [1:0] MP1_9_out_demux_peripheral_mscbus;
wire            MP2_0_IO;
wire      [4:0] MP2_0_in_mux_en_mscbus;
wire      [4:0] MP2_0_in_mux_peripheral_mscbus;
wire      [2:0] MP2_0_out_demux_peripheral_mscbus;
wire            MP2_10_IO;
wire      [3:0] MP2_10_in_mux_en_mscbus;
wire      [3:0] MP2_10_in_mux_peripheral_mscbus;
wire      [1:0] MP2_10_out_demux_peripheral_mscbus;
wire            MP2_11_IO;
wire      [2:0] MP2_11_in_mux_en_mscbus;
wire      [2:0] MP2_11_in_mux_peripheral_mscbus;
wire      [2:0] MP2_11_out_demux_peripheral_mscbus;
wire            MP2_12_IO;
wire      [2:0] MP2_12_in_mux_en_mscbus;
wire      [2:0] MP2_12_in_mux_peripheral_mscbus;
wire      [2:0] MP2_12_out_demux_peripheral_mscbus;
wire            MP2_13_IO;
wire      [1:0] MP2_13_in_mux_en_mscbus;
wire      [1:0] MP2_13_in_mux_peripheral_mscbus;
wire      [3:0] MP2_13_out_demux_peripheral_mscbus;
wire            MP2_14_IO;
wire      [3:0] MP2_14_in_mux_en_mscbus;
wire      [3:0] MP2_14_in_mux_peripheral_mscbus;
wire      [1:0] MP2_14_out_demux_peripheral_mscbus;
wire            MP2_15_IO;
wire      [1:0] MP2_15_in_mux_en_mscbus;
wire      [1:0] MP2_15_in_mux_peripheral_mscbus;
wire      [3:0] MP2_15_out_demux_peripheral_mscbus;
wire            MP2_1_IO;
wire      [2:0] MP2_1_in_mux_en_mscbus;
wire      [2:0] MP2_1_in_mux_peripheral_mscbus;
wire      [4:0] MP2_1_out_demux_peripheral_mscbus;
wire            MP2_2_IO;
wire      [4:0] MP2_2_in_mux_en_mscbus;
wire      [4:0] MP2_2_in_mux_peripheral_mscbus;
wire      [2:0] MP2_2_out_demux_peripheral_mscbus;
wire            MP2_3_IO;
wire      [3:0] MP2_3_in_mux_en_mscbus;
wire      [3:0] MP2_3_in_mux_peripheral_mscbus;
wire      [3:0] MP2_3_out_demux_peripheral_mscbus;
wire            MP2_4_IO;
wire      [4:0] MP2_4_in_mux_en_mscbus;
wire      [4:0] MP2_4_in_mux_peripheral_mscbus;
wire      [2:0] MP2_4_out_demux_peripheral_mscbus;
wire            MP2_5_IO;
wire      [3:0] MP2_5_in_mux_en_mscbus;
wire      [3:0] MP2_5_in_mux_peripheral_mscbus;
wire      [3:0] MP2_5_out_demux_peripheral_mscbus;
wire            MP2_6_IO;
wire      [4:0] MP2_6_in_mux_en_mscbus;
wire      [4:0] MP2_6_in_mux_peripheral_mscbus;
wire      [2:0] MP2_6_out_demux_peripheral_mscbus;
wire            MP2_7_IO;
wire      [3:0] MP2_7_in_mux_en_mscbus;
wire      [3:0] MP2_7_in_mux_peripheral_mscbus;
wire      [3:0] MP2_7_out_demux_peripheral_mscbus;
wire            MP2_8_IO;
wire      [2:0] MP2_8_in_mux_en_mscbus;
wire      [2:0] MP2_8_in_mux_peripheral_mscbus;
wire      [1:0] MP2_8_out_demux_peripheral_mscbus;
wire            MP2_9_IO;
wire      [1:0] MP2_9_in_mux_en_mscbus;
wire      [1:0] MP2_9_in_mux_peripheral_mscbus;
wire      [3:0] MP2_9_out_demux_peripheral_mscbus;
wire            PWR_ON_RSTn_IO;
wire            RESETOUTn_IO;
wire            SGMII0RXN_IO;
wire            SGMII0RXP_IO;
wire            SGMII0TXN_IO;
wire            SGMII0TXP_IO;
wire            SGMII1RXN_IO;
wire            SGMII1RXP_IO;
wire            SGMII1TXN_IO;
wire            SGMII1TXP_IO;
wire            SGMII2RXN_IO;
wire            SGMII2RXP_IO;
wire            SGMII2TXN_IO;
wire            SGMII2TXP_IO;
wire            SPI0LPBCLKUNB_IO;
wire            SPI1LPBCLKUNB_IO;
wire            SPI2LPBCLKUNB_IO;
wire            SPI3LPBCLKUNB_IO;
wire            SPI4LPBCLKUNB_IO;
wire            SPI5LPBCLKUNB_IO;
wire            SPI6LPBCLKUNB_IO;
wire            SPI7LPBCLKUNB_IO;
wire            SPI8LPBCLKUNB_IO;
wire            SPI9LPBCLKUNB_IO;
wire            TCK_IO;
wire            TDI_IO;
wire            TDO_IO;
wire            TMS_IO;
wire            TRSTN_IO;
wire            VDDS_REF0_HI_IO;
wire            VDDS_REF0_LO_IO;
wire            VDDS_REF1_HI_IO;
wire            VDDS_REF1_LO_IO;
wire            VDDS_REF2_HI_IO;
wire            VDDS_REF2_LO_IO;
wire            VDDS_REF_LPD_HI_IO;
wire            VDDS_REF_LPD_LO_IO;
wire            VDDS_REF_SD_HI_IO;
wire            VDDS_REF_SD_LO_IO;
wire            X1_IO;
wire            X2_IO;
wire            XSPI0LBCLKUNB_IO;
wire            gpio_clock;
wire            gpio_reset_n;
wire            io_ADC0EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC0EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC0EXTMUXSEL0_adcchsel;
wire            io_ADC0EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC0EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC0EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC0EXTMUXSEL0_adcofftrim;
wire            io_ADC0EXTMUXSEL0_adcpwrdn;
wire            io_ADC0EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC0EXTMUXSEL0_adcresult;
wire            io_ADC0EXTMUXSEL0_adcsignalmode;
wire            io_ADC0EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC0EXTMUXSEL0_dtb;
wire            io_ADC0EXTMUXSEL0_samcapreset_disable;
wire            io_ADC0EXTMUXSEL0_samcapreset_level;
wire            io_ADC0EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC0EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC0EXTMUXSEL1_adcchsel;
wire            io_ADC0EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC0EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC0EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC0EXTMUXSEL1_adcofftrim;
wire            io_ADC0EXTMUXSEL1_adcpwrdn;
wire            io_ADC0EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC0EXTMUXSEL1_adcresult;
wire            io_ADC0EXTMUXSEL1_adcsignalmode;
wire            io_ADC0EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC0EXTMUXSEL1_dtb;
wire            io_ADC0EXTMUXSEL1_samcapreset_disable;
wire            io_ADC0EXTMUXSEL1_samcapreset_level;
wire            io_ADC0EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC0EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC0EXTMUXSEL2_adcchsel;
wire            io_ADC0EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC0EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC0EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC0EXTMUXSEL2_adcofftrim;
wire            io_ADC0EXTMUXSEL2_adcpwrdn;
wire            io_ADC0EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC0EXTMUXSEL2_adcresult;
wire            io_ADC0EXTMUXSEL2_adcsignalmode;
wire            io_ADC0EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC0EXTMUXSEL2_dtb;
wire            io_ADC0EXTMUXSEL2_samcapreset_disable;
wire            io_ADC0EXTMUXSEL2_samcapreset_level;
wire            io_ADC0EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC0EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC0EXTMUXSEL3_adcchsel;
wire            io_ADC0EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC0EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC0EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC0EXTMUXSEL3_adcofftrim;
wire            io_ADC0EXTMUXSEL3_adcpwrdn;
wire            io_ADC0EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC0EXTMUXSEL3_adcresult;
wire            io_ADC0EXTMUXSEL3_adcsignalmode;
wire            io_ADC0EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC0EXTMUXSEL3_dtb;
wire            io_ADC0EXTMUXSEL3_samcapreset_disable;
wire            io_ADC0EXTMUXSEL3_samcapreset_level;
wire            io_ADC1EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC1EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC1EXTMUXSEL0_adcchsel;
wire            io_ADC1EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC1EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC1EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC1EXTMUXSEL0_adcofftrim;
wire            io_ADC1EXTMUXSEL0_adcpwrdn;
wire            io_ADC1EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC1EXTMUXSEL0_adcresult;
wire            io_ADC1EXTMUXSEL0_adcsignalmode;
wire            io_ADC1EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC1EXTMUXSEL0_dtb;
wire            io_ADC1EXTMUXSEL0_samcapreset_disable;
wire            io_ADC1EXTMUXSEL0_samcapreset_level;
wire            io_ADC1EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC1EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC1EXTMUXSEL1_adcchsel;
wire            io_ADC1EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC1EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC1EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC1EXTMUXSEL1_adcofftrim;
wire            io_ADC1EXTMUXSEL1_adcpwrdn;
wire            io_ADC1EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC1EXTMUXSEL1_adcresult;
wire            io_ADC1EXTMUXSEL1_adcsignalmode;
wire            io_ADC1EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC1EXTMUXSEL1_dtb;
wire            io_ADC1EXTMUXSEL1_samcapreset_disable;
wire            io_ADC1EXTMUXSEL1_samcapreset_level;
wire            io_ADC1EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC1EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC1EXTMUXSEL2_adcchsel;
wire            io_ADC1EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC1EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC1EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC1EXTMUXSEL2_adcofftrim;
wire            io_ADC1EXTMUXSEL2_adcpwrdn;
wire            io_ADC1EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC1EXTMUXSEL2_adcresult;
wire            io_ADC1EXTMUXSEL2_adcsignalmode;
wire            io_ADC1EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC1EXTMUXSEL2_dtb;
wire            io_ADC1EXTMUXSEL2_samcapreset_disable;
wire            io_ADC1EXTMUXSEL2_samcapreset_level;
wire            io_ADC1EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC1EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC1EXTMUXSEL3_adcchsel;
wire            io_ADC1EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC1EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC1EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC1EXTMUXSEL3_adcofftrim;
wire            io_ADC1EXTMUXSEL3_adcpwrdn;
wire            io_ADC1EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC1EXTMUXSEL3_adcresult;
wire            io_ADC1EXTMUXSEL3_adcsignalmode;
wire            io_ADC1EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC1EXTMUXSEL3_dtb;
wire            io_ADC1EXTMUXSEL3_samcapreset_disable;
wire            io_ADC1EXTMUXSEL3_samcapreset_level;
wire            io_ADC2EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC2EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC2EXTMUXSEL0_adcchsel;
wire            io_ADC2EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC2EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC2EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC2EXTMUXSEL0_adcofftrim;
wire            io_ADC2EXTMUXSEL0_adcpwrdn;
wire            io_ADC2EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC2EXTMUXSEL0_adcresult;
wire            io_ADC2EXTMUXSEL0_adcsignalmode;
wire            io_ADC2EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC2EXTMUXSEL0_dtb;
wire            io_ADC2EXTMUXSEL0_samcapreset_disable;
wire            io_ADC2EXTMUXSEL0_samcapreset_level;
wire            io_ADC2EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC2EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC2EXTMUXSEL1_adcchsel;
wire            io_ADC2EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC2EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC2EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC2EXTMUXSEL1_adcofftrim;
wire            io_ADC2EXTMUXSEL1_adcpwrdn;
wire            io_ADC2EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC2EXTMUXSEL1_adcresult;
wire            io_ADC2EXTMUXSEL1_adcsignalmode;
wire            io_ADC2EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC2EXTMUXSEL1_dtb;
wire            io_ADC2EXTMUXSEL1_samcapreset_disable;
wire            io_ADC2EXTMUXSEL1_samcapreset_level;
wire            io_ADC2EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC2EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC2EXTMUXSEL2_adcchsel;
wire            io_ADC2EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC2EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC2EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC2EXTMUXSEL2_adcofftrim;
wire            io_ADC2EXTMUXSEL2_adcpwrdn;
wire            io_ADC2EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC2EXTMUXSEL2_adcresult;
wire            io_ADC2EXTMUXSEL2_adcsignalmode;
wire            io_ADC2EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC2EXTMUXSEL2_dtb;
wire            io_ADC2EXTMUXSEL2_samcapreset_disable;
wire            io_ADC2EXTMUXSEL2_samcapreset_level;
wire            io_ADC2EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC2EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC2EXTMUXSEL3_adcchsel;
wire            io_ADC2EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC2EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC2EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC2EXTMUXSEL3_adcofftrim;
wire            io_ADC2EXTMUXSEL3_adcpwrdn;
wire            io_ADC2EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC2EXTMUXSEL3_adcresult;
wire            io_ADC2EXTMUXSEL3_adcsignalmode;
wire            io_ADC2EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC2EXTMUXSEL3_dtb;
wire            io_ADC2EXTMUXSEL3_samcapreset_disable;
wire            io_ADC2EXTMUXSEL3_samcapreset_level;
wire            io_ADC3EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC3EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC3EXTMUXSEL0_adcchsel;
wire            io_ADC3EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC3EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC3EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC3EXTMUXSEL0_adcofftrim;
wire            io_ADC3EXTMUXSEL0_adcpwrdn;
wire            io_ADC3EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC3EXTMUXSEL0_adcresult;
wire            io_ADC3EXTMUXSEL0_adcsignalmode;
wire            io_ADC3EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC3EXTMUXSEL0_dtb;
wire            io_ADC3EXTMUXSEL0_samcapreset_disable;
wire            io_ADC3EXTMUXSEL0_samcapreset_level;
wire            io_ADC3EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC3EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC3EXTMUXSEL1_adcchsel;
wire            io_ADC3EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC3EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC3EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC3EXTMUXSEL1_adcofftrim;
wire            io_ADC3EXTMUXSEL1_adcpwrdn;
wire            io_ADC3EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC3EXTMUXSEL1_adcresult;
wire            io_ADC3EXTMUXSEL1_adcsignalmode;
wire            io_ADC3EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC3EXTMUXSEL1_dtb;
wire            io_ADC3EXTMUXSEL1_samcapreset_disable;
wire            io_ADC3EXTMUXSEL1_samcapreset_level;
wire            io_ADC3EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC3EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC3EXTMUXSEL2_adcchsel;
wire            io_ADC3EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC3EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC3EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC3EXTMUXSEL2_adcofftrim;
wire            io_ADC3EXTMUXSEL2_adcpwrdn;
wire            io_ADC3EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC3EXTMUXSEL2_adcresult;
wire            io_ADC3EXTMUXSEL2_adcsignalmode;
wire            io_ADC3EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC3EXTMUXSEL2_dtb;
wire            io_ADC3EXTMUXSEL2_samcapreset_disable;
wire            io_ADC3EXTMUXSEL2_samcapreset_level;
wire            io_ADC3EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC3EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC3EXTMUXSEL3_adcchsel;
wire            io_ADC3EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC3EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC3EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC3EXTMUXSEL3_adcofftrim;
wire            io_ADC3EXTMUXSEL3_adcpwrdn;
wire            io_ADC3EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC3EXTMUXSEL3_adcresult;
wire            io_ADC3EXTMUXSEL3_adcsignalmode;
wire            io_ADC3EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC3EXTMUXSEL3_dtb;
wire            io_ADC3EXTMUXSEL3_samcapreset_disable;
wire            io_ADC3EXTMUXSEL3_samcapreset_level;
wire            io_ADC4EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC4EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC4EXTMUXSEL0_adcchsel;
wire            io_ADC4EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC4EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC4EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC4EXTMUXSEL0_adcofftrim;
wire            io_ADC4EXTMUXSEL0_adcpwrdn;
wire            io_ADC4EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC4EXTMUXSEL0_adcresult;
wire            io_ADC4EXTMUXSEL0_adcsignalmode;
wire            io_ADC4EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC4EXTMUXSEL0_dtb;
wire            io_ADC4EXTMUXSEL0_samcapreset_disable;
wire            io_ADC4EXTMUXSEL0_samcapreset_level;
wire            io_ADC4EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC4EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC4EXTMUXSEL1_adcchsel;
wire            io_ADC4EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC4EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC4EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC4EXTMUXSEL1_adcofftrim;
wire            io_ADC4EXTMUXSEL1_adcpwrdn;
wire            io_ADC4EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC4EXTMUXSEL1_adcresult;
wire            io_ADC4EXTMUXSEL1_adcsignalmode;
wire            io_ADC4EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC4EXTMUXSEL1_dtb;
wire            io_ADC4EXTMUXSEL1_samcapreset_disable;
wire            io_ADC4EXTMUXSEL1_samcapreset_level;
wire            io_ADC4EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC4EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC4EXTMUXSEL2_adcchsel;
wire            io_ADC4EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC4EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC4EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC4EXTMUXSEL2_adcofftrim;
wire            io_ADC4EXTMUXSEL2_adcpwrdn;
wire            io_ADC4EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC4EXTMUXSEL2_adcresult;
wire            io_ADC4EXTMUXSEL2_adcsignalmode;
wire            io_ADC4EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC4EXTMUXSEL2_dtb;
wire            io_ADC4EXTMUXSEL2_samcapreset_disable;
wire            io_ADC4EXTMUXSEL2_samcapreset_level;
wire            io_ADC4EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC4EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC4EXTMUXSEL3_adcchsel;
wire            io_ADC4EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC4EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC4EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC4EXTMUXSEL3_adcofftrim;
wire            io_ADC4EXTMUXSEL3_adcpwrdn;
wire            io_ADC4EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC4EXTMUXSEL3_adcresult;
wire            io_ADC4EXTMUXSEL3_adcsignalmode;
wire            io_ADC4EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC4EXTMUXSEL3_dtb;
wire            io_ADC4EXTMUXSEL3_samcapreset_disable;
wire            io_ADC4EXTMUXSEL3_samcapreset_level;
wire            io_ADC5EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC5EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC5EXTMUXSEL0_adcchsel;
wire            io_ADC5EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC5EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC5EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC5EXTMUXSEL0_adcofftrim;
wire            io_ADC5EXTMUXSEL0_adcpwrdn;
wire            io_ADC5EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC5EXTMUXSEL0_adcresult;
wire            io_ADC5EXTMUXSEL0_adcsignalmode;
wire            io_ADC5EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC5EXTMUXSEL0_dtb;
wire            io_ADC5EXTMUXSEL0_samcapreset_disable;
wire            io_ADC5EXTMUXSEL0_samcapreset_level;
wire            io_ADC5EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC5EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC5EXTMUXSEL1_adcchsel;
wire            io_ADC5EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC5EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC5EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC5EXTMUXSEL1_adcofftrim;
wire            io_ADC5EXTMUXSEL1_adcpwrdn;
wire            io_ADC5EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC5EXTMUXSEL1_adcresult;
wire            io_ADC5EXTMUXSEL1_adcsignalmode;
wire            io_ADC5EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC5EXTMUXSEL1_dtb;
wire            io_ADC5EXTMUXSEL1_samcapreset_disable;
wire            io_ADC5EXTMUXSEL1_samcapreset_level;
wire            io_ADC5EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC5EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC5EXTMUXSEL2_adcchsel;
wire            io_ADC5EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC5EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC5EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC5EXTMUXSEL2_adcofftrim;
wire            io_ADC5EXTMUXSEL2_adcpwrdn;
wire            io_ADC5EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC5EXTMUXSEL2_adcresult;
wire            io_ADC5EXTMUXSEL2_adcsignalmode;
wire            io_ADC5EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC5EXTMUXSEL2_dtb;
wire            io_ADC5EXTMUXSEL2_samcapreset_disable;
wire            io_ADC5EXTMUXSEL2_samcapreset_level;
wire            io_ADC5EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC5EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC5EXTMUXSEL3_adcchsel;
wire            io_ADC5EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC5EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC5EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC5EXTMUXSEL3_adcofftrim;
wire            io_ADC5EXTMUXSEL3_adcpwrdn;
wire            io_ADC5EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC5EXTMUXSEL3_adcresult;
wire            io_ADC5EXTMUXSEL3_adcsignalmode;
wire            io_ADC5EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC5EXTMUXSEL3_dtb;
wire            io_ADC5EXTMUXSEL3_samcapreset_disable;
wire            io_ADC5EXTMUXSEL3_samcapreset_level;
wire            io_ADC6EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC6EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC6EXTMUXSEL0_adcchsel;
wire            io_ADC6EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC6EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC6EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC6EXTMUXSEL0_adcofftrim;
wire            io_ADC6EXTMUXSEL0_adcpwrdn;
wire            io_ADC6EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC6EXTMUXSEL0_adcresult;
wire            io_ADC6EXTMUXSEL0_adcsignalmode;
wire            io_ADC6EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC6EXTMUXSEL0_dtb;
wire            io_ADC6EXTMUXSEL0_samcapreset_disable;
wire            io_ADC6EXTMUXSEL0_samcapreset_level;
wire            io_ADC6EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC6EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC6EXTMUXSEL1_adcchsel;
wire            io_ADC6EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC6EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC6EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC6EXTMUXSEL1_adcofftrim;
wire            io_ADC6EXTMUXSEL1_adcpwrdn;
wire            io_ADC6EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC6EXTMUXSEL1_adcresult;
wire            io_ADC6EXTMUXSEL1_adcsignalmode;
wire            io_ADC6EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC6EXTMUXSEL1_dtb;
wire            io_ADC6EXTMUXSEL1_samcapreset_disable;
wire            io_ADC6EXTMUXSEL1_samcapreset_level;
wire            io_ADC6EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC6EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC6EXTMUXSEL2_adcchsel;
wire            io_ADC6EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC6EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC6EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC6EXTMUXSEL2_adcofftrim;
wire            io_ADC6EXTMUXSEL2_adcpwrdn;
wire            io_ADC6EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC6EXTMUXSEL2_adcresult;
wire            io_ADC6EXTMUXSEL2_adcsignalmode;
wire            io_ADC6EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC6EXTMUXSEL2_dtb;
wire            io_ADC6EXTMUXSEL2_samcapreset_disable;
wire            io_ADC6EXTMUXSEL2_samcapreset_level;
wire            io_ADC6EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC6EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC6EXTMUXSEL3_adcchsel;
wire            io_ADC6EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC6EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC6EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC6EXTMUXSEL3_adcofftrim;
wire            io_ADC6EXTMUXSEL3_adcpwrdn;
wire            io_ADC6EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC6EXTMUXSEL3_adcresult;
wire            io_ADC6EXTMUXSEL3_adcsignalmode;
wire            io_ADC6EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC6EXTMUXSEL3_dtb;
wire            io_ADC6EXTMUXSEL3_samcapreset_disable;
wire            io_ADC6EXTMUXSEL3_samcapreset_level;
wire            io_ADC7EXTMUXSEL0_adccalibmode;
wire      [4:0] io_ADC7EXTMUXSEL0_adccalibstep;
wire      [4:0] io_ADC7EXTMUXSEL0_adcchsel;
wire            io_ADC7EXTMUXSEL0_adcclk;
wire     [31:0] io_ADC7EXTMUXSEL0_adcconfig;
wire     [31:0] io_ADC7EXTMUXSEL0_adcinltrim1;
wire     [15:0] io_ADC7EXTMUXSEL0_adcofftrim;
wire            io_ADC7EXTMUXSEL0_adcpwrdn;
wire            io_ADC7EXTMUXSEL0_adcresolution;
wire     [15:0] io_ADC7EXTMUXSEL0_adcresult;
wire            io_ADC7EXTMUXSEL0_adcsignalmode;
wire            io_ADC7EXTMUXSEL0_adcsoc;
wire     [15:0] io_ADC7EXTMUXSEL0_dtb;
wire            io_ADC7EXTMUXSEL0_samcapreset_disable;
wire            io_ADC7EXTMUXSEL0_samcapreset_level;
wire            io_ADC7EXTMUXSEL1_adccalibmode;
wire      [4:0] io_ADC7EXTMUXSEL1_adccalibstep;
wire      [4:0] io_ADC7EXTMUXSEL1_adcchsel;
wire            io_ADC7EXTMUXSEL1_adcclk;
wire     [31:0] io_ADC7EXTMUXSEL1_adcconfig;
wire     [31:0] io_ADC7EXTMUXSEL1_adcinltrim1;
wire     [15:0] io_ADC7EXTMUXSEL1_adcofftrim;
wire            io_ADC7EXTMUXSEL1_adcpwrdn;
wire            io_ADC7EXTMUXSEL1_adcresolution;
wire     [15:0] io_ADC7EXTMUXSEL1_adcresult;
wire            io_ADC7EXTMUXSEL1_adcsignalmode;
wire            io_ADC7EXTMUXSEL1_adcsoc;
wire     [15:0] io_ADC7EXTMUXSEL1_dtb;
wire            io_ADC7EXTMUXSEL1_samcapreset_disable;
wire            io_ADC7EXTMUXSEL1_samcapreset_level;
wire            io_ADC7EXTMUXSEL2_adccalibmode;
wire      [4:0] io_ADC7EXTMUXSEL2_adccalibstep;
wire      [4:0] io_ADC7EXTMUXSEL2_adcchsel;
wire            io_ADC7EXTMUXSEL2_adcclk;
wire     [31:0] io_ADC7EXTMUXSEL2_adcconfig;
wire     [31:0] io_ADC7EXTMUXSEL2_adcinltrim1;
wire     [15:0] io_ADC7EXTMUXSEL2_adcofftrim;
wire            io_ADC7EXTMUXSEL2_adcpwrdn;
wire            io_ADC7EXTMUXSEL2_adcresolution;
wire     [15:0] io_ADC7EXTMUXSEL2_adcresult;
wire            io_ADC7EXTMUXSEL2_adcsignalmode;
wire            io_ADC7EXTMUXSEL2_adcsoc;
wire     [15:0] io_ADC7EXTMUXSEL2_dtb;
wire            io_ADC7EXTMUXSEL2_samcapreset_disable;
wire            io_ADC7EXTMUXSEL2_samcapreset_level;
wire            io_ADC7EXTMUXSEL3_adccalibmode;
wire      [4:0] io_ADC7EXTMUXSEL3_adccalibstep;
wire      [4:0] io_ADC7EXTMUXSEL3_adcchsel;
wire            io_ADC7EXTMUXSEL3_adcclk;
wire     [31:0] io_ADC7EXTMUXSEL3_adcconfig;
wire     [31:0] io_ADC7EXTMUXSEL3_adcinltrim1;
wire     [15:0] io_ADC7EXTMUXSEL3_adcofftrim;
wire            io_ADC7EXTMUXSEL3_adcpwrdn;
wire            io_ADC7EXTMUXSEL3_adcresolution;
wire     [15:0] io_ADC7EXTMUXSEL3_adcresult;
wire            io_ADC7EXTMUXSEL3_adcsignalmode;
wire            io_ADC7EXTMUXSEL3_adcsoc;
wire     [15:0] io_ADC7EXTMUXSEL3_dtb;
wire            io_ADC7EXTMUXSEL3_samcapreset_disable;
wire            io_ADC7EXTMUXSEL3_samcapreset_level;
wire            io_ADCSOC0_adccalibmode;
wire      [4:0] io_ADCSOC0_adccalibstep;
wire      [4:0] io_ADCSOC0_adcchsel;
wire            io_ADCSOC0_adcclk;
wire     [31:0] io_ADCSOC0_adcconfig;
wire     [31:0] io_ADCSOC0_adcinltrim1;
wire     [15:0] io_ADCSOC0_adcofftrim;
wire            io_ADCSOC0_adcpwrdn;
wire            io_ADCSOC0_adcresolution;
wire     [15:0] io_ADCSOC0_adcresult;
wire            io_ADCSOC0_adcsignalmode;
wire            io_ADCSOC0_adcsoc;
wire     [15:0] io_ADCSOC0_dtb;
wire            io_ADCSOC0_samcapreset_disable;
wire            io_ADCSOC0_samcapreset_level;
wire            io_ADCSOC1_adccalibmode;
wire      [4:0] io_ADCSOC1_adccalibstep;
wire      [4:0] io_ADCSOC1_adcchsel;
wire            io_ADCSOC1_adcclk;
wire     [31:0] io_ADCSOC1_adcconfig;
wire     [31:0] io_ADCSOC1_adcinltrim1;
wire     [15:0] io_ADCSOC1_adcofftrim;
wire            io_ADCSOC1_adcpwrdn;
wire            io_ADCSOC1_adcresolution;
wire     [15:0] io_ADCSOC1_adcresult;
wire            io_ADCSOC1_adcsignalmode;
wire            io_ADCSOC1_adcsoc;
wire     [15:0] io_ADCSOC1_dtb;
wire            io_ADCSOC1_samcapreset_disable;
wire            io_ADCSOC1_samcapreset_level;
wire            io_CAN0_rxd;
wire            io_CAN0_txd;
wire            io_CAN10_rxd;
wire            io_CAN10_txd;
wire            io_CAN11_rxd;
wire            io_CAN11_txd;
wire            io_CAN1_rxd;
wire            io_CAN1_txd;
wire            io_CAN2_rxd;
wire            io_CAN2_txd;
wire            io_CAN3_rxd;
wire            io_CAN3_txd;
wire            io_CAN4_rxd;
wire            io_CAN4_txd;
wire            io_CAN5_rxd;
wire            io_CAN5_txd;
wire            io_CAN6_rxd;
wire            io_CAN6_txd;
wire            io_CAN7_rxd;
wire            io_CAN7_txd;
wire            io_CAN8_rxd;
wire            io_CAN8_txd;
wire            io_CAN9_rxd;
wire            io_CAN9_txd;
wire            io_EPWM0_a_i;
wire            io_EPWM0_a_o;
wire            io_EPWM0_a_oen;
wire            io_EPWM0_b_i;
wire            io_EPWM0_b_o;
wire            io_EPWM0_b_oen;
wire            io_EPWM10_a_i;
wire            io_EPWM10_a_o;
wire            io_EPWM10_a_oen;
wire            io_EPWM10_b_i;
wire            io_EPWM10_b_o;
wire            io_EPWM10_b_oen;
wire            io_EPWM11_a_i;
wire            io_EPWM11_a_o;
wire            io_EPWM11_a_oen;
wire            io_EPWM11_b_i;
wire            io_EPWM11_b_o;
wire            io_EPWM11_b_oen;
wire            io_EPWM12_a_i;
wire            io_EPWM12_a_o;
wire            io_EPWM12_a_oen;
wire            io_EPWM12_b_i;
wire            io_EPWM12_b_o;
wire            io_EPWM12_b_oen;
wire            io_EPWM13_a_i;
wire            io_EPWM13_a_o;
wire            io_EPWM13_a_oen;
wire            io_EPWM13_b_i;
wire            io_EPWM13_b_o;
wire            io_EPWM13_b_oen;
wire            io_EPWM14_a_i;
wire            io_EPWM14_a_o;
wire            io_EPWM14_a_oen;
wire            io_EPWM14_b_i;
wire            io_EPWM14_b_o;
wire            io_EPWM14_b_oen;
wire            io_EPWM15_a_i;
wire            io_EPWM15_a_o;
wire            io_EPWM15_a_oen;
wire            io_EPWM15_b_i;
wire            io_EPWM15_b_o;
wire            io_EPWM15_b_oen;
wire            io_EPWM16_a_i;
wire            io_EPWM16_a_o;
wire            io_EPWM16_a_oen;
wire            io_EPWM16_b_i;
wire            io_EPWM16_b_o;
wire            io_EPWM16_b_oen;
wire            io_EPWM17_a_i;
wire            io_EPWM17_a_o;
wire            io_EPWM17_a_oen;
wire            io_EPWM17_b_i;
wire            io_EPWM17_b_o;
wire            io_EPWM17_b_oen;
wire            io_EPWM18_a_i;
wire            io_EPWM18_a_o;
wire            io_EPWM18_a_oen;
wire            io_EPWM18_b_i;
wire            io_EPWM18_b_o;
wire            io_EPWM18_b_oen;
wire            io_EPWM19_a_i;
wire            io_EPWM19_a_o;
wire            io_EPWM19_a_oen;
wire            io_EPWM19_b_i;
wire            io_EPWM19_b_o;
wire            io_EPWM19_b_oen;
wire            io_EPWM1_a_i;
wire            io_EPWM1_a_o;
wire            io_EPWM1_a_oen;
wire            io_EPWM1_b_i;
wire            io_EPWM1_b_o;
wire            io_EPWM1_b_oen;
wire            io_EPWM20_a_i;
wire            io_EPWM20_a_o;
wire            io_EPWM20_a_oen;
wire            io_EPWM20_b_i;
wire            io_EPWM20_b_o;
wire            io_EPWM20_b_oen;
wire            io_EPWM21_a_i;
wire            io_EPWM21_a_o;
wire            io_EPWM21_a_oen;
wire            io_EPWM21_b_i;
wire            io_EPWM21_b_o;
wire            io_EPWM21_b_oen;
wire            io_EPWM22_a_i;
wire            io_EPWM22_a_o;
wire            io_EPWM22_a_oen;
wire            io_EPWM22_b_i;
wire            io_EPWM22_b_o;
wire            io_EPWM22_b_oen;
wire            io_EPWM23_a_i;
wire            io_EPWM23_a_o;
wire            io_EPWM23_a_oen;
wire            io_EPWM23_b_i;
wire            io_EPWM23_b_o;
wire            io_EPWM23_b_oen;
wire            io_EPWM24_a_i;
wire            io_EPWM24_a_o;
wire            io_EPWM24_a_oen;
wire            io_EPWM24_b_i;
wire            io_EPWM24_b_o;
wire            io_EPWM24_b_oen;
wire            io_EPWM25_a_i;
wire            io_EPWM25_a_o;
wire            io_EPWM25_a_oen;
wire            io_EPWM25_b_i;
wire            io_EPWM25_b_o;
wire            io_EPWM25_b_oen;
wire            io_EPWM26_a_i;
wire            io_EPWM26_a_o;
wire            io_EPWM26_a_oen;
wire            io_EPWM26_b_i;
wire            io_EPWM26_b_o;
wire            io_EPWM26_b_oen;
wire            io_EPWM27_a_i;
wire            io_EPWM27_a_o;
wire            io_EPWM27_a_oen;
wire            io_EPWM27_b_i;
wire            io_EPWM27_b_o;
wire            io_EPWM27_b_oen;
wire            io_EPWM28_a_i;
wire            io_EPWM28_a_o;
wire            io_EPWM28_a_oen;
wire            io_EPWM28_b_i;
wire            io_EPWM28_b_o;
wire            io_EPWM28_b_oen;
wire            io_EPWM29_a_i;
wire            io_EPWM29_a_o;
wire            io_EPWM29_a_oen;
wire            io_EPWM29_b_i;
wire            io_EPWM29_b_o;
wire            io_EPWM29_b_oen;
wire            io_EPWM2_a_i;
wire            io_EPWM2_a_o;
wire            io_EPWM2_a_oen;
wire            io_EPWM2_b_i;
wire            io_EPWM2_b_o;
wire            io_EPWM2_b_oen;
wire            io_EPWM30_a_i;
wire            io_EPWM30_a_o;
wire            io_EPWM30_a_oen;
wire            io_EPWM30_b_i;
wire            io_EPWM30_b_o;
wire            io_EPWM30_b_oen;
wire            io_EPWM31_a_i;
wire            io_EPWM31_a_o;
wire            io_EPWM31_a_oen;
wire            io_EPWM31_b_i;
wire            io_EPWM31_b_o;
wire            io_EPWM31_b_oen;
wire            io_EPWM3_a_i;
wire            io_EPWM3_a_o;
wire            io_EPWM3_a_oen;
wire            io_EPWM3_b_i;
wire            io_EPWM3_b_o;
wire            io_EPWM3_b_oen;
wire            io_EPWM4_a_i;
wire            io_EPWM4_a_o;
wire            io_EPWM4_a_oen;
wire            io_EPWM4_b_i;
wire            io_EPWM4_b_o;
wire            io_EPWM4_b_oen;
wire            io_EPWM5_a_i;
wire            io_EPWM5_a_o;
wire            io_EPWM5_a_oen;
wire            io_EPWM5_b_i;
wire            io_EPWM5_b_o;
wire            io_EPWM5_b_oen;
wire            io_EPWM6_a_i;
wire            io_EPWM6_a_o;
wire            io_EPWM6_a_oen;
wire            io_EPWM6_b_i;
wire            io_EPWM6_b_o;
wire            io_EPWM6_b_oen;
wire            io_EPWM7_a_i;
wire            io_EPWM7_a_o;
wire            io_EPWM7_a_oen;
wire            io_EPWM7_b_i;
wire            io_EPWM7_b_o;
wire            io_EPWM7_b_oen;
wire            io_EPWM8_a_i;
wire            io_EPWM8_a_o;
wire            io_EPWM8_a_oen;
wire            io_EPWM8_b_i;
wire            io_EPWM8_b_o;
wire            io_EPWM8_b_oen;
wire            io_EPWM9_a_i;
wire            io_EPWM9_a_o;
wire            io_EPWM9_a_oen;
wire            io_EPWM9_b_i;
wire            io_EPWM9_b_o;
wire            io_EPWM9_b_oen;
wire            io_EPWMSYNCO_a_i;
wire            io_EPWMSYNCO_a_o;
wire            io_EPWMSYNCO_a_oen;
wire            io_EPWMSYNCO_b_i;
wire            io_EPWMSYNCO_b_o;
wire            io_EPWMSYNCO_b_oen;
wire            io_FSI0RX_ck;
wire            io_FSI0RX_d0;
wire            io_FSI0RX_d1;
wire            io_FSI0TX_ck;
wire            io_FSI0TX_d0;
wire            io_FSI0TX_d1;
wire            io_FSI1RX_ck;
wire            io_FSI1RX_d0;
wire            io_FSI1RX_d1;
wire            io_FSI1TX_ck;
wire            io_FSI1TX_d0;
wire            io_FSI1TX_d1;
wire            io_FSI2RX_ck;
wire            io_FSI2RX_d0;
wire            io_FSI2RX_d1;
wire            io_FSI2TX_ck;
wire            io_FSI2TX_d0;
wire            io_FSI2TX_d1;
wire            io_FSI3RX_ck;
wire            io_FSI3RX_d0;
wire            io_FSI3RX_d1;
wire            io_FSI3TX_ck;
wire            io_FSI3TX_d0;
wire            io_FSI3TX_d1;
wire            io_FSI4RX_ck;
wire            io_FSI4RX_d0;
wire            io_FSI4RX_d1;
wire            io_FSI4TX_ck;
wire            io_FSI4TX_d0;
wire            io_FSI4TX_d1;
wire            io_FSI5RX_ck;
wire            io_FSI5RX_d0;
wire            io_FSI5RX_d1;
wire            io_FSI5TX_ck;
wire            io_FSI5TX_d0;
wire            io_FSI5TX_d1;
wire            io_I2C0SCL_piscl;
wire            io_I2C0SCL_pisda;
wire            io_I2C0SCL_porsccbe;
wire            io_I2C0SCL_porscl;
wire            io_I2C0SCL_porsclhsmode;
wire            io_I2C0SCL_porsclnmode;
wire            io_I2C0SCL_porsda;
wire            io_I2C0SCL_porsdagzn;
wire            io_I2C0SCL_porsdanmode;
wire            io_I2C0SCL_porsdhsmode;
wire            io_I2C1SCL_piscl;
wire            io_I2C1SCL_pisda;
wire            io_I2C1SCL_porsccbe;
wire            io_I2C1SCL_porscl;
wire            io_I2C1SCL_porsclhsmode;
wire            io_I2C1SCL_porsclnmode;
wire            io_I2C1SCL_porsda;
wire            io_I2C1SCL_porsdagzn;
wire            io_I2C1SCL_porsdanmode;
wire            io_I2C1SCL_porsdhsmode;
wire            io_I2C2SCL_piscl;
wire            io_I2C2SCL_pisda;
wire            io_I2C2SCL_porsccbe;
wire            io_I2C2SCL_porscl;
wire            io_I2C2SCL_porsclhsmode;
wire            io_I2C2SCL_porsclnmode;
wire            io_I2C2SCL_porsda;
wire            io_I2C2SCL_porsdagzn;
wire            io_I2C2SCL_porsdanmode;
wire            io_I2C2SCL_porsdhsmode;
wire            io_I2C3SCL_piscl;
wire            io_I2C3SCL_pisda;
wire            io_I2C3SCL_porsccbe;
wire            io_I2C3SCL_porscl;
wire            io_I2C3SCL_porsclhsmode;
wire            io_I2C3SCL_porsclnmode;
wire            io_I2C3SCL_porsda;
wire            io_I2C3SCL_porsdagzn;
wire            io_I2C3SCL_porsdanmode;
wire            io_I2C3SCL_porsdhsmode;
wire            io_LIN0_rxd;
wire            io_LIN0_tr_en;
wire            io_LIN0_txd;
wire            io_LIN1_rxd;
wire            io_LIN1_tr_en;
wire            io_LIN1_txd;
wire            io_LIN2_rxd;
wire            io_LIN2_tr_en;
wire            io_LIN2_txd;
wire            io_LIN3_rxd;
wire            io_LIN3_tr_en;
wire            io_LIN3_txd;
wire            io_LIN4_rxd;
wire            io_LIN4_tr_en;
wire            io_LIN4_txd;
wire            io_LIN5_rxd;
wire            io_LIN5_tr_en;
wire            io_LIN5_txd;
wire            io_LIN6_rxd;
wire            io_LIN6_tr_en;
wire            io_LIN6_txd;
wire            io_LIN7_rxd;
wire            io_LIN7_tr_en;
wire            io_LIN7_txd;
wire            io_LPD_CAN0RX_rxd;
wire            io_LPD_CAN0RX_txd;
wire            io_LPD_CAN0TX_rxd;
wire            io_LPD_CAN0TX_txd;
wire            io_LPD_LIN0RX_rxd;
wire            io_LPD_LIN0RX_tr_en;
wire            io_LPD_LIN0RX_txd;
wire            io_LPD_LIN0TX_rxd;
wire            io_LPD_LIN0TX_tr_en;
wire            io_LPD_LIN0TX_txd;
wire            io_MIBSPI0CLK_clock;
wire            io_MIBSPI0CS0_in;
wire            io_MIBSPI0CS0_oen;
wire            io_MIBSPI0CS0_out;
wire            io_MIBSPI0CS10_in;
wire            io_MIBSPI0CS10_oen;
wire            io_MIBSPI0CS10_out;
wire            io_MIBSPI0CS11_in;
wire            io_MIBSPI0CS11_oen;
wire            io_MIBSPI0CS11_out;
wire            io_MIBSPI0CS1_in;
wire            io_MIBSPI0CS1_oen;
wire            io_MIBSPI0CS1_out;
wire            io_MIBSPI0CS2_in;
wire            io_MIBSPI0CS2_oen;
wire            io_MIBSPI0CS2_out;
wire            io_MIBSPI0CS3_in;
wire            io_MIBSPI0CS3_oen;
wire            io_MIBSPI0CS3_out;
wire            io_MIBSPI0CS4_in;
wire            io_MIBSPI0CS4_oen;
wire            io_MIBSPI0CS4_out;
wire            io_MIBSPI0CS5_in;
wire            io_MIBSPI0CS5_oen;
wire            io_MIBSPI0CS5_out;
wire            io_MIBSPI0CS6_in;
wire            io_MIBSPI0CS6_oen;
wire            io_MIBSPI0CS6_out;
wire            io_MIBSPI0CS7_in;
wire            io_MIBSPI0CS7_oen;
wire            io_MIBSPI0CS7_out;
wire            io_MIBSPI0CS8_in;
wire            io_MIBSPI0CS8_oen;
wire            io_MIBSPI0CS8_out;
wire            io_MIBSPI0CS9_in;
wire            io_MIBSPI0CS9_oen;
wire            io_MIBSPI0CS9_out;
wire            io_MIBSPI0PICO_in;
wire            io_MIBSPI0PICO_oen;
wire            io_MIBSPI0PICO_out;
wire            io_MIBSPI0POCI_in;
wire            io_MIBSPI0POCI_oen;
wire            io_MIBSPI0POCI_out;
wire            io_MIBSPI1CLK_clock;
wire            io_MIBSPI1CS0_in;
wire            io_MIBSPI1CS0_oen;
wire            io_MIBSPI1CS0_out;
wire            io_MIBSPI1CS10_in;
wire            io_MIBSPI1CS10_oen;
wire            io_MIBSPI1CS10_out;
wire            io_MIBSPI1CS11_in;
wire            io_MIBSPI1CS11_oen;
wire            io_MIBSPI1CS11_out;
wire            io_MIBSPI1CS1_in;
wire            io_MIBSPI1CS1_oen;
wire            io_MIBSPI1CS1_out;
wire            io_MIBSPI1CS2_in;
wire            io_MIBSPI1CS2_oen;
wire            io_MIBSPI1CS2_out;
wire            io_MIBSPI1CS3_in;
wire            io_MIBSPI1CS3_oen;
wire            io_MIBSPI1CS3_out;
wire            io_MIBSPI1CS4_in;
wire            io_MIBSPI1CS4_oen;
wire            io_MIBSPI1CS4_out;
wire            io_MIBSPI1CS5_in;
wire            io_MIBSPI1CS5_oen;
wire            io_MIBSPI1CS5_out;
wire            io_MIBSPI1CS6_in;
wire            io_MIBSPI1CS6_oen;
wire            io_MIBSPI1CS6_out;
wire            io_MIBSPI1CS7_in;
wire            io_MIBSPI1CS7_oen;
wire            io_MIBSPI1CS7_out;
wire            io_MIBSPI1CS8_in;
wire            io_MIBSPI1CS8_oen;
wire            io_MIBSPI1CS8_out;
wire            io_MIBSPI1CS9_in;
wire            io_MIBSPI1CS9_oen;
wire            io_MIBSPI1CS9_out;
wire            io_MIBSPI1PICO_in;
wire            io_MIBSPI1PICO_oen;
wire            io_MIBSPI1PICO_out;
wire            io_MIBSPI1POCI_in;
wire            io_MIBSPI1POCI_oen;
wire            io_MIBSPI1POCI_out;
wire            io_OUTPUTXBAR0_intr;
wire            io_OUTPUTXBAR10_intr;
wire            io_OUTPUTXBAR11_intr;
wire            io_OUTPUTXBAR12_intr;
wire            io_OUTPUTXBAR13_intr;
wire            io_OUTPUTXBAR14_intr;
wire            io_OUTPUTXBAR15_intr;
wire            io_OUTPUTXBAR1_intr;
wire            io_OUTPUTXBAR2_intr;
wire            io_OUTPUTXBAR3_intr;
wire            io_OUTPUTXBAR4_intr;
wire            io_OUTPUTXBAR5_intr;
wire            io_OUTPUTXBAR6_intr;
wire            io_OUTPUTXBAR7_intr;
wire            io_OUTPUTXBAR8_intr;
wire            io_OUTPUTXBAR9_intr;
wire      [3:0] io_PSI5_0_rx;
wire      [3:0] io_PSI5_0_tx;
wire      [3:0] io_PSI5_1_rx;
wire      [3:0] io_PSI5_1_tx;
wire      [3:0] io_PSI5_2_rx;
wire      [3:0] io_PSI5_2_tx;
wire      [3:0] io_PSI5_3_rx;
wire      [3:0] io_PSI5_3_tx;
wire            io_SDFM0_i_clock1;
wire            io_SDFM0_i_clock2;
wire            io_SDFM0_i_clock3;
wire            io_SDFM0_i_clock4;
wire            io_SDFM0_i_datain1;
wire            io_SDFM0_i_datain2;
wire            io_SDFM0_i_datain3;
wire            io_SDFM0_i_datain4;
wire            io_SDFM10_i_clock1;
wire            io_SDFM10_i_clock2;
wire            io_SDFM10_i_clock3;
wire            io_SDFM10_i_clock4;
wire            io_SDFM10_i_datain1;
wire            io_SDFM10_i_datain2;
wire            io_SDFM10_i_datain3;
wire            io_SDFM10_i_datain4;
wire            io_SDFM11_i_clock1;
wire            io_SDFM11_i_clock2;
wire            io_SDFM11_i_clock3;
wire            io_SDFM11_i_clock4;
wire            io_SDFM11_i_datain1;
wire            io_SDFM11_i_datain2;
wire            io_SDFM11_i_datain3;
wire            io_SDFM11_i_datain4;
wire            io_SDFM1_i_clock1;
wire            io_SDFM1_i_clock2;
wire            io_SDFM1_i_clock3;
wire            io_SDFM1_i_clock4;
wire            io_SDFM1_i_datain1;
wire            io_SDFM1_i_datain2;
wire            io_SDFM1_i_datain3;
wire            io_SDFM1_i_datain4;
wire            io_SDFM2_i_clock1;
wire            io_SDFM2_i_clock2;
wire            io_SDFM2_i_clock3;
wire            io_SDFM2_i_clock4;
wire            io_SDFM2_i_datain1;
wire            io_SDFM2_i_datain2;
wire            io_SDFM2_i_datain3;
wire            io_SDFM2_i_datain4;
wire            io_SDFM3_i_clock1;
wire            io_SDFM3_i_clock2;
wire            io_SDFM3_i_clock3;
wire            io_SDFM3_i_clock4;
wire            io_SDFM3_i_datain1;
wire            io_SDFM3_i_datain2;
wire            io_SDFM3_i_datain3;
wire            io_SDFM3_i_datain4;
wire            io_SDFM4_i_clock1;
wire            io_SDFM4_i_clock2;
wire            io_SDFM4_i_clock3;
wire            io_SDFM4_i_clock4;
wire            io_SDFM4_i_datain1;
wire            io_SDFM4_i_datain2;
wire            io_SDFM4_i_datain3;
wire            io_SDFM4_i_datain4;
wire            io_SDFM5_i_clock1;
wire            io_SDFM5_i_clock2;
wire            io_SDFM5_i_clock3;
wire            io_SDFM5_i_clock4;
wire            io_SDFM5_i_datain1;
wire            io_SDFM5_i_datain2;
wire            io_SDFM5_i_datain3;
wire            io_SDFM5_i_datain4;
wire            io_SDFM6_i_clock1;
wire            io_SDFM6_i_clock2;
wire            io_SDFM6_i_clock3;
wire            io_SDFM6_i_clock4;
wire            io_SDFM6_i_datain1;
wire            io_SDFM6_i_datain2;
wire            io_SDFM6_i_datain3;
wire            io_SDFM6_i_datain4;
wire            io_SDFM7_i_clock1;
wire            io_SDFM7_i_clock2;
wire            io_SDFM7_i_clock3;
wire            io_SDFM7_i_clock4;
wire            io_SDFM7_i_datain1;
wire            io_SDFM7_i_datain2;
wire            io_SDFM7_i_datain3;
wire            io_SDFM7_i_datain4;
wire            io_SDFM8_i_clock1;
wire            io_SDFM8_i_clock2;
wire            io_SDFM8_i_clock3;
wire            io_SDFM8_i_clock4;
wire            io_SDFM8_i_datain1;
wire            io_SDFM8_i_datain2;
wire            io_SDFM8_i_datain3;
wire            io_SDFM8_i_datain4;
wire            io_SDFM9_i_clock1;
wire            io_SDFM9_i_clock2;
wire            io_SDFM9_i_clock3;
wire            io_SDFM9_i_clock4;
wire            io_SDFM9_i_datain1;
wire            io_SDFM9_i_datain2;
wire            io_SDFM9_i_datain3;
wire            io_SDFM9_i_datain4;
wire            io_SENT0_rxd_i;
wire            io_SENT0_rxd_o;
wire            io_SENT0_rxd_oen_o;
wire    [121:0] io_SENT0_soc_ext_trig_i;
wire     [31:0] io_SENT0_tstamp_val_i;
wire            io_SENT1_rxd_i;
wire            io_SENT1_rxd_o;
wire            io_SENT1_rxd_oen_o;
wire    [121:0] io_SENT1_soc_ext_trig_i;
wire     [31:0] io_SENT1_tstamp_val_i;
wire            io_SENT2_rxd_i;
wire            io_SENT2_rxd_o;
wire            io_SENT2_rxd_oen_o;
wire    [121:0] io_SENT2_soc_ext_trig_i;
wire     [31:0] io_SENT2_tstamp_val_i;
wire            io_SENT3_rxd_i;
wire            io_SENT3_rxd_o;
wire            io_SENT3_rxd_oen_o;
wire    [121:0] io_SENT3_soc_ext_trig_i;
wire     [31:0] io_SENT3_tstamp_val_i;
wire            io_SENT4_rxd_i;
wire            io_SENT4_rxd_o;
wire            io_SENT4_rxd_oen_o;
wire    [121:0] io_SENT4_soc_ext_trig_i;
wire     [31:0] io_SENT4_tstamp_val_i;
wire            io_SENT5_rxd_i;
wire            io_SENT5_rxd_o;
wire            io_SENT5_rxd_oen_o;
wire    [121:0] io_SENT5_soc_ext_trig_i;
wire     [31:0] io_SENT5_tstamp_val_i;
wire            io_SPI2CLK_clock;
wire            io_SPI2CS0_in;
wire            io_SPI2CS0_oen;
wire            io_SPI2CS0_out;
wire            io_SPI2CS1_in;
wire            io_SPI2CS1_oen;
wire            io_SPI2CS1_out;
wire            io_SPI2CS2_in;
wire            io_SPI2CS2_oen;
wire            io_SPI2CS2_out;
wire            io_SPI2CS3_in;
wire            io_SPI2CS3_oen;
wire            io_SPI2CS3_out;
wire            io_SPI2CS4_in;
wire            io_SPI2CS4_oen;
wire            io_SPI2CS4_out;
wire            io_SPI2CS5_in;
wire            io_SPI2CS5_oen;
wire            io_SPI2CS5_out;
wire            io_SPI2PICO_in;
wire            io_SPI2PICO_oen;
wire            io_SPI2PICO_out;
wire            io_SPI2POCI_in;
wire            io_SPI2POCI_oen;
wire            io_SPI2POCI_out;
wire            io_SPI3CLK_clock;
wire            io_SPI3CS0_in;
wire            io_SPI3CS0_oen;
wire            io_SPI3CS0_out;
wire            io_SPI3CS1_in;
wire            io_SPI3CS1_oen;
wire            io_SPI3CS1_out;
wire            io_SPI3CS2_in;
wire            io_SPI3CS2_oen;
wire            io_SPI3CS2_out;
wire            io_SPI3CS3_in;
wire            io_SPI3CS3_oen;
wire            io_SPI3CS3_out;
wire            io_SPI3CS4_in;
wire            io_SPI3CS4_oen;
wire            io_SPI3CS4_out;
wire            io_SPI3CS5_in;
wire            io_SPI3CS5_oen;
wire            io_SPI3CS5_out;
wire            io_SPI3PICO_in;
wire            io_SPI3PICO_oen;
wire            io_SPI3PICO_out;
wire            io_SPI3POCI_in;
wire            io_SPI3POCI_oen;
wire            io_SPI3POCI_out;
wire            io_SPI4CLK_clock;
wire            io_SPI4CS0_in;
wire            io_SPI4CS0_oen;
wire            io_SPI4CS0_out;
wire            io_SPI4CS1_in;
wire            io_SPI4CS1_oen;
wire            io_SPI4CS1_out;
wire            io_SPI4CS2_in;
wire            io_SPI4CS2_oen;
wire            io_SPI4CS2_out;
wire            io_SPI4CS3_in;
wire            io_SPI4CS3_oen;
wire            io_SPI4CS3_out;
wire            io_SPI4CS4_in;
wire            io_SPI4CS4_oen;
wire            io_SPI4CS4_out;
wire            io_SPI4CS5_in;
wire            io_SPI4CS5_oen;
wire            io_SPI4CS5_out;
wire            io_SPI4PICO_in;
wire            io_SPI4PICO_oen;
wire            io_SPI4PICO_out;
wire            io_SPI4POCI_in;
wire            io_SPI4POCI_oen;
wire            io_SPI4POCI_out;
wire            io_SPI5CLK_clock;
wire            io_SPI5CS0_in;
wire            io_SPI5CS0_oen;
wire            io_SPI5CS0_out;
wire            io_SPI5CS1_in;
wire            io_SPI5CS1_oen;
wire            io_SPI5CS1_out;
wire            io_SPI5CS2_in;
wire            io_SPI5CS2_oen;
wire            io_SPI5CS2_out;
wire            io_SPI5CS3_in;
wire            io_SPI5CS3_oen;
wire            io_SPI5CS3_out;
wire            io_SPI5CS4_in;
wire            io_SPI5CS4_oen;
wire            io_SPI5CS4_out;
wire            io_SPI5CS5_in;
wire            io_SPI5CS5_oen;
wire            io_SPI5CS5_out;
wire            io_SPI5PICO_in;
wire            io_SPI5PICO_oen;
wire            io_SPI5PICO_out;
wire            io_SPI5POCI_in;
wire            io_SPI5POCI_oen;
wire            io_SPI5POCI_out;
wire            io_SPI6CLK_clock;
wire            io_SPI6CS0_in;
wire            io_SPI6CS0_oen;
wire            io_SPI6CS0_out;
wire            io_SPI6CS1_in;
wire            io_SPI6CS1_oen;
wire            io_SPI6CS1_out;
wire            io_SPI6CS2_in;
wire            io_SPI6CS2_oen;
wire            io_SPI6CS2_out;
wire            io_SPI6CS3_in;
wire            io_SPI6CS3_oen;
wire            io_SPI6CS3_out;
wire            io_SPI6CS4_in;
wire            io_SPI6CS4_oen;
wire            io_SPI6CS4_out;
wire            io_SPI6CS5_in;
wire            io_SPI6CS5_oen;
wire            io_SPI6CS5_out;
wire            io_SPI6PICO_in;
wire            io_SPI6PICO_oen;
wire            io_SPI6PICO_out;
wire            io_SPI6POCI_in;
wire            io_SPI6POCI_oen;
wire            io_SPI6POCI_out;
wire            io_SPI7CLK_clock;
wire            io_SPI7CS0_in;
wire            io_SPI7CS0_oen;
wire            io_SPI7CS0_out;
wire            io_SPI7CS1_in;
wire            io_SPI7CS1_oen;
wire            io_SPI7CS1_out;
wire            io_SPI7CS2_in;
wire            io_SPI7CS2_oen;
wire            io_SPI7CS2_out;
wire            io_SPI7CS3_in;
wire            io_SPI7CS3_oen;
wire            io_SPI7CS3_out;
wire            io_SPI7CS4_in;
wire            io_SPI7CS4_oen;
wire            io_SPI7CS4_out;
wire            io_SPI7CS5_in;
wire            io_SPI7CS5_oen;
wire            io_SPI7CS5_out;
wire            io_SPI7PICO_in;
wire            io_SPI7PICO_oen;
wire            io_SPI7PICO_out;
wire            io_SPI7POCI_in;
wire            io_SPI7POCI_oen;
wire            io_SPI7POCI_out;
wire            io_SPI8CLK_clock;
wire            io_SPI8CS0_in;
wire            io_SPI8CS0_oen;
wire            io_SPI8CS0_out;
wire            io_SPI8CS1_in;
wire            io_SPI8CS1_oen;
wire            io_SPI8CS1_out;
wire            io_SPI8CS2_in;
wire            io_SPI8CS2_oen;
wire            io_SPI8CS2_out;
wire            io_SPI8CS3_in;
wire            io_SPI8CS3_oen;
wire            io_SPI8CS3_out;
wire            io_SPI8CS4_in;
wire            io_SPI8CS4_oen;
wire            io_SPI8CS4_out;
wire            io_SPI8CS5_in;
wire            io_SPI8CS5_oen;
wire            io_SPI8CS5_out;
wire            io_SPI8PICO_in;
wire            io_SPI8PICO_oen;
wire            io_SPI8PICO_out;
wire            io_SPI8POCI_in;
wire            io_SPI8POCI_oen;
wire            io_SPI8POCI_out;
wire            io_SPI9CLK_clock;
wire            io_SPI9CS0_in;
wire            io_SPI9CS0_oen;
wire            io_SPI9CS0_out;
wire            io_SPI9CS1_in;
wire            io_SPI9CS1_oen;
wire            io_SPI9CS1_out;
wire            io_SPI9CS2_in;
wire            io_SPI9CS2_oen;
wire            io_SPI9CS2_out;
wire            io_SPI9CS3_in;
wire            io_SPI9CS3_oen;
wire            io_SPI9CS3_out;
wire            io_SPI9CS4_in;
wire            io_SPI9CS4_oen;
wire            io_SPI9CS4_out;
wire            io_SPI9CS5_in;
wire            io_SPI9CS5_oen;
wire            io_SPI9CS5_out;
wire            io_SPI9PICO_in;
wire            io_SPI9PICO_oen;
wire            io_SPI9PICO_out;
wire            io_SPI9POCI_in;
wire            io_SPI9POCI_oen;
wire            io_SPI9POCI_out;
wire            io_UART0_cd_n;
wire            io_UART0_cts_n;
wire            io_UART0_dsr_n;
wire            io_UART0_dtr_n;
wire            io_UART0_out1;
wire            io_UART0_out2;
wire            io_UART0_ri_n;
wire            io_UART0_rts_n;
wire            io_UART0_rx;
wire            io_UART0_tx;
wire            io_UART1_cd_n;
wire            io_UART1_cts_n;
wire            io_UART1_dsr_n;
wire            io_UART1_dtr_n;
wire            io_UART1_out1;
wire            io_UART1_out2;
wire            io_UART1_ri_n;
wire            io_UART1_rts_n;
wire            io_UART1_rx;
wire            io_UART1_tx;
wire      [3:0] io_XSPI0_cs_o;
wire      [7:0] io_XSPI0_data_i;
wire            io_XSPI0_data_mask_o;
wire            io_XSPI0_data_mask_oe_n;
wire      [7:0] io_XSPI0_data_o;
wire      [7:0] io_XSPI0_data_oe_n;
wire            io_XSPI0_dqs_clk;
wire      [3:0] io_XSPI0_intr_n;
wire            io_XSPI0_mst_in_clk;
wire            io_XSPI0_out_clk;
wire      [3:0] io_XSPI0_reset_in;
wire      [3:0] io_XSPI0_reset_out;
wire     [31:0] io_ap0_GP_DATA_IN_out_mscbus;
wire     [31:0] io_ap0_amsel_out_mscbus;
wire     [31:0] io_ap0_async_in_from_pad_mscbus;
wire     [31:0] io_ap0_data_out_2_pinmux_mscbus;
wire     [31:0] io_ap0_dir_out_mscbus;
wire     [31:0] io_ap0_ds0_out_mscbus;
wire     [31:0] io_ap0_ds1_out_mscbus;
wire     [31:0] io_ap0_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_ap0_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_ap0_gpio_out_2_buf_mscbus;
wire     [31:0] io_ap0_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_ap0_in_function_en_out_mscbus;
wire     [31:0] io_ap0_in_termination_en_out_mscbus;
wire     [31:0] io_ap0_inena_out_mscbus;
wire     [31:0] io_ap0_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_ap0_mode0_out_mscbus;
wire     [31:0] io_ap0_mode1_out_mscbus;
wire    [255:0] io_ap0_pes_en_out_mscbus;
wire     [31:0] io_ap0_pes_in_en_out_mscbus;
wire     [63:0] io_ap0_pes_safeval_out_mscbus;
wire    [159:0] io_ap0_pinmux_muxsel_out_mscbus;
wire     [31:0] io_ap0_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_ap0_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_ap0_pull_en_out_mscbus;
wire     [31:0] io_ap0_pull_type_out_mscbus;
wire     [31:0] io_ap0_schmitt_out_mscbus;
wire     [31:0] io_ap0_slew_out_mscbus;
wire     [31:0] io_ap1_GP_DATA_IN_out_mscbus;
wire     [31:0] io_ap1_amsel_out_mscbus;
wire     [31:0] io_ap1_async_in_from_pad_mscbus;
wire     [31:0] io_ap1_data_out_2_pinmux_mscbus;
wire     [31:0] io_ap1_dir_out_mscbus;
wire     [31:0] io_ap1_ds0_out_mscbus;
wire     [31:0] io_ap1_ds1_out_mscbus;
wire     [31:0] io_ap1_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_ap1_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_ap1_gpio_out_2_buf_mscbus;
wire     [31:0] io_ap1_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_ap1_in_function_en_out_mscbus;
wire     [31:0] io_ap1_in_termination_en_out_mscbus;
wire     [31:0] io_ap1_inena_out_mscbus;
wire     [31:0] io_ap1_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_ap1_mode0_out_mscbus;
wire     [31:0] io_ap1_mode1_out_mscbus;
wire    [255:0] io_ap1_pes_en_out_mscbus;
wire     [31:0] io_ap1_pes_in_en_out_mscbus;
wire     [63:0] io_ap1_pes_safeval_out_mscbus;
wire    [159:0] io_ap1_pinmux_muxsel_out_mscbus;
wire     [31:0] io_ap1_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_ap1_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_ap1_pull_en_out_mscbus;
wire     [31:0] io_ap1_pull_type_out_mscbus;
wire     [31:0] io_ap1_schmitt_out_mscbus;
wire     [31:0] io_ap1_slew_out_mscbus;
wire            io_clock;
wire     [31:0] io_dp0_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp0_amsel_out_mscbus;
wire     [31:0] io_dp0_async_in_from_pad_mscbus;
wire     [31:0] io_dp0_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp0_dir_out_mscbus;
wire     [31:0] io_dp0_ds0_out_mscbus;
wire     [31:0] io_dp0_ds1_out_mscbus;
wire     [31:0] io_dp0_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp0_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp0_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp0_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp0_in_function_en_out_mscbus;
wire     [31:0] io_dp0_in_termination_en_out_mscbus;
wire     [31:0] io_dp0_inena_out_mscbus;
wire     [31:0] io_dp0_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp0_mode0_out_mscbus;
wire     [31:0] io_dp0_mode1_out_mscbus;
wire    [255:0] io_dp0_pes_en_out_mscbus;
wire     [31:0] io_dp0_pes_in_en_out_mscbus;
wire     [63:0] io_dp0_pes_safeval_out_mscbus;
wire    [159:0] io_dp0_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp0_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp0_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp0_pull_en_out_mscbus;
wire     [31:0] io_dp0_pull_type_out_mscbus;
wire     [31:0] io_dp0_schmitt_out_mscbus;
wire     [31:0] io_dp0_slew_out_mscbus;
wire     [31:0] io_dp1_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp1_amsel_out_mscbus;
wire     [31:0] io_dp1_async_in_from_pad_mscbus;
wire     [31:0] io_dp1_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp1_dir_out_mscbus;
wire     [31:0] io_dp1_ds0_out_mscbus;
wire     [31:0] io_dp1_ds1_out_mscbus;
wire     [31:0] io_dp1_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp1_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp1_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp1_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp1_in_function_en_out_mscbus;
wire     [31:0] io_dp1_in_termination_en_out_mscbus;
wire     [31:0] io_dp1_inena_out_mscbus;
wire     [31:0] io_dp1_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp1_mode0_out_mscbus;
wire     [31:0] io_dp1_mode1_out_mscbus;
wire    [255:0] io_dp1_pes_en_out_mscbus;
wire     [31:0] io_dp1_pes_in_en_out_mscbus;
wire     [63:0] io_dp1_pes_safeval_out_mscbus;
wire    [159:0] io_dp1_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp1_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp1_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp1_pull_en_out_mscbus;
wire     [31:0] io_dp1_pull_type_out_mscbus;
wire     [31:0] io_dp1_schmitt_out_mscbus;
wire     [31:0] io_dp1_slew_out_mscbus;
wire     [31:0] io_dp2_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp2_amsel_out_mscbus;
wire     [31:0] io_dp2_async_in_from_pad_mscbus;
wire     [31:0] io_dp2_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp2_dir_out_mscbus;
wire     [31:0] io_dp2_ds0_out_mscbus;
wire     [31:0] io_dp2_ds1_out_mscbus;
wire     [31:0] io_dp2_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp2_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp2_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp2_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp2_in_function_en_out_mscbus;
wire     [31:0] io_dp2_in_termination_en_out_mscbus;
wire     [31:0] io_dp2_inena_out_mscbus;
wire     [31:0] io_dp2_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp2_mode0_out_mscbus;
wire     [31:0] io_dp2_mode1_out_mscbus;
wire    [255:0] io_dp2_pes_en_out_mscbus;
wire     [31:0] io_dp2_pes_in_en_out_mscbus;
wire     [63:0] io_dp2_pes_safeval_out_mscbus;
wire    [159:0] io_dp2_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp2_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp2_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp2_pull_en_out_mscbus;
wire     [31:0] io_dp2_pull_type_out_mscbus;
wire     [31:0] io_dp2_schmitt_out_mscbus;
wire     [31:0] io_dp2_slew_out_mscbus;
wire     [31:0] io_dp3_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp3_amsel_out_mscbus;
wire     [31:0] io_dp3_async_in_from_pad_mscbus;
wire     [31:0] io_dp3_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp3_dir_out_mscbus;
wire     [31:0] io_dp3_ds0_out_mscbus;
wire     [31:0] io_dp3_ds1_out_mscbus;
wire     [31:0] io_dp3_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp3_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp3_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp3_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp3_in_function_en_out_mscbus;
wire     [31:0] io_dp3_in_termination_en_out_mscbus;
wire     [31:0] io_dp3_inena_out_mscbus;
wire     [31:0] io_dp3_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp3_mode0_out_mscbus;
wire     [31:0] io_dp3_mode1_out_mscbus;
wire    [255:0] io_dp3_pes_en_out_mscbus;
wire     [31:0] io_dp3_pes_in_en_out_mscbus;
wire     [63:0] io_dp3_pes_safeval_out_mscbus;
wire    [159:0] io_dp3_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp3_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp3_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp3_pull_en_out_mscbus;
wire     [31:0] io_dp3_pull_type_out_mscbus;
wire     [31:0] io_dp3_schmitt_out_mscbus;
wire     [31:0] io_dp3_slew_out_mscbus;
wire     [31:0] io_dp4_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp4_amsel_out_mscbus;
wire     [31:0] io_dp4_async_in_from_pad_mscbus;
wire     [31:0] io_dp4_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp4_dir_out_mscbus;
wire     [31:0] io_dp4_ds0_out_mscbus;
wire     [31:0] io_dp4_ds1_out_mscbus;
wire     [31:0] io_dp4_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp4_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp4_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp4_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp4_in_function_en_out_mscbus;
wire     [31:0] io_dp4_in_termination_en_out_mscbus;
wire     [31:0] io_dp4_inena_out_mscbus;
wire     [31:0] io_dp4_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp4_mode0_out_mscbus;
wire     [31:0] io_dp4_mode1_out_mscbus;
wire    [255:0] io_dp4_pes_en_out_mscbus;
wire     [31:0] io_dp4_pes_in_en_out_mscbus;
wire     [63:0] io_dp4_pes_safeval_out_mscbus;
wire    [159:0] io_dp4_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp4_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp4_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp4_pull_en_out_mscbus;
wire     [31:0] io_dp4_pull_type_out_mscbus;
wire     [31:0] io_dp4_schmitt_out_mscbus;
wire     [31:0] io_dp4_slew_out_mscbus;
wire     [31:0] io_dp5_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp5_amsel_out_mscbus;
wire     [31:0] io_dp5_async_in_from_pad_mscbus;
wire     [31:0] io_dp5_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp5_dir_out_mscbus;
wire     [31:0] io_dp5_ds0_out_mscbus;
wire     [31:0] io_dp5_ds1_out_mscbus;
wire     [31:0] io_dp5_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp5_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp5_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp5_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp5_in_function_en_out_mscbus;
wire     [31:0] io_dp5_in_termination_en_out_mscbus;
wire     [31:0] io_dp5_inena_out_mscbus;
wire     [31:0] io_dp5_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp5_mode0_out_mscbus;
wire     [31:0] io_dp5_mode1_out_mscbus;
wire    [255:0] io_dp5_pes_en_out_mscbus;
wire     [31:0] io_dp5_pes_in_en_out_mscbus;
wire     [63:0] io_dp5_pes_safeval_out_mscbus;
wire    [159:0] io_dp5_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp5_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp5_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp5_pull_en_out_mscbus;
wire     [31:0] io_dp5_pull_type_out_mscbus;
wire     [31:0] io_dp5_schmitt_out_mscbus;
wire     [31:0] io_dp5_slew_out_mscbus;
wire     [31:0] io_dp6_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp6_amsel_out_mscbus;
wire     [31:0] io_dp6_async_in_from_pad_mscbus;
wire     [31:0] io_dp6_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp6_dir_out_mscbus;
wire     [31:0] io_dp6_ds0_out_mscbus;
wire     [31:0] io_dp6_ds1_out_mscbus;
wire     [31:0] io_dp6_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp6_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp6_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp6_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp6_in_function_en_out_mscbus;
wire     [31:0] io_dp6_in_termination_en_out_mscbus;
wire     [31:0] io_dp6_inena_out_mscbus;
wire     [31:0] io_dp6_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp6_mode0_out_mscbus;
wire     [31:0] io_dp6_mode1_out_mscbus;
wire    [255:0] io_dp6_pes_en_out_mscbus;
wire     [31:0] io_dp6_pes_in_en_out_mscbus;
wire     [63:0] io_dp6_pes_safeval_out_mscbus;
wire    [159:0] io_dp6_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp6_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp6_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp6_pull_en_out_mscbus;
wire     [31:0] io_dp6_pull_type_out_mscbus;
wire     [31:0] io_dp6_schmitt_out_mscbus;
wire     [31:0] io_dp6_slew_out_mscbus;
wire     [31:0] io_dp7_GP_DATA_IN_out_mscbus;
wire     [31:0] io_dp7_amsel_out_mscbus;
wire     [31:0] io_dp7_async_in_from_pad_mscbus;
wire     [31:0] io_dp7_data_out_2_pinmux_mscbus;
wire     [31:0] io_dp7_dir_out_mscbus;
wire     [31:0] io_dp7_ds0_out_mscbus;
wire     [31:0] io_dp7_ds1_out_mscbus;
wire     [31:0] io_dp7_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_dp7_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_dp7_gpio_out_2_buf_mscbus;
wire     [31:0] io_dp7_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_dp7_in_function_en_out_mscbus;
wire     [31:0] io_dp7_in_termination_en_out_mscbus;
wire     [31:0] io_dp7_inena_out_mscbus;
wire     [31:0] io_dp7_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_dp7_mode0_out_mscbus;
wire     [31:0] io_dp7_mode1_out_mscbus;
wire    [255:0] io_dp7_pes_en_out_mscbus;
wire     [31:0] io_dp7_pes_in_en_out_mscbus;
wire     [63:0] io_dp7_pes_safeval_out_mscbus;
wire    [159:0] io_dp7_pinmux_muxsel_out_mscbus;
wire     [31:0] io_dp7_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_dp7_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_dp7_pull_en_out_mscbus;
wire     [31:0] io_dp7_pull_type_out_mscbus;
wire     [31:0] io_dp7_schmitt_out_mscbus;
wire     [31:0] io_dp7_slew_out_mscbus;
wire      [4:0] io_ext_ADC0EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC0EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC0EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC0EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC1EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC1EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC1EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC1EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC2EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC2EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC2EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC2EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC3EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC3EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC3EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC3EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC4EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC4EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC4EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC4EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC5EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC5EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC5EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC5EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC6EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC6EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC6EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC6EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADC7EXTMUXSEL0_adcchsel;
wire      [4:0] io_ext_ADC7EXTMUXSEL1_adcchsel;
wire      [4:0] io_ext_ADC7EXTMUXSEL2_adcchsel;
wire      [4:0] io_ext_ADC7EXTMUXSEL3_adcchsel;
wire      [4:0] io_ext_ADCSOC0_adcchsel;
wire      [4:0] io_ext_ADCSOC1_adcchsel;
wire     [31:0] io_mp0_GP_DATA_IN_out_mscbus;
wire     [31:0] io_mp0_amsel_out_mscbus;
wire     [31:0] io_mp0_async_in_from_pad_mscbus;
wire     [31:0] io_mp0_data_out_2_pinmux_mscbus;
wire     [31:0] io_mp0_dir_out_mscbus;
wire     [31:0] io_mp0_ds0_out_mscbus;
wire     [31:0] io_mp0_ds1_out_mscbus;
wire     [31:0] io_mp0_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_mp0_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_mp0_gpio_out_2_buf_mscbus;
wire     [31:0] io_mp0_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_mp0_in_function_en_out_mscbus;
wire     [31:0] io_mp0_in_termination_en_out_mscbus;
wire     [31:0] io_mp0_inena_out_mscbus;
wire     [31:0] io_mp0_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_mp0_mode0_out_mscbus;
wire     [31:0] io_mp0_mode1_out_mscbus;
wire    [255:0] io_mp0_pes_en_out_mscbus;
wire     [31:0] io_mp0_pes_in_en_out_mscbus;
wire     [63:0] io_mp0_pes_safeval_out_mscbus;
wire    [159:0] io_mp0_pinmux_muxsel_out_mscbus;
wire     [31:0] io_mp0_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_mp0_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_mp0_pull_en_out_mscbus;
wire     [31:0] io_mp0_pull_type_out_mscbus;
wire     [31:0] io_mp0_schmitt_out_mscbus;
wire     [31:0] io_mp0_slew_out_mscbus;
wire     [31:0] io_mp1_GP_DATA_IN_out_mscbus;
wire     [31:0] io_mp1_amsel_out_mscbus;
wire     [31:0] io_mp1_async_in_from_pad_mscbus;
wire     [31:0] io_mp1_data_out_2_pinmux_mscbus;
wire     [31:0] io_mp1_dir_out_mscbus;
wire     [31:0] io_mp1_ds0_out_mscbus;
wire     [31:0] io_mp1_ds1_out_mscbus;
wire     [31:0] io_mp1_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_mp1_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_mp1_gpio_out_2_buf_mscbus;
wire     [31:0] io_mp1_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_mp1_in_function_en_out_mscbus;
wire     [31:0] io_mp1_in_termination_en_out_mscbus;
wire     [31:0] io_mp1_inena_out_mscbus;
wire     [31:0] io_mp1_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_mp1_mode0_out_mscbus;
wire     [31:0] io_mp1_mode1_out_mscbus;
wire    [255:0] io_mp1_pes_en_out_mscbus;
wire     [31:0] io_mp1_pes_in_en_out_mscbus;
wire     [63:0] io_mp1_pes_safeval_out_mscbus;
wire    [159:0] io_mp1_pinmux_muxsel_out_mscbus;
wire     [31:0] io_mp1_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_mp1_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_mp1_pull_en_out_mscbus;
wire     [31:0] io_mp1_pull_type_out_mscbus;
wire     [31:0] io_mp1_schmitt_out_mscbus;
wire     [31:0] io_mp1_slew_out_mscbus;
wire     [31:0] io_mp2_GP_DATA_IN_out_mscbus;
wire     [31:0] io_mp2_amsel_out_mscbus;
wire     [31:0] io_mp2_async_in_from_pad_mscbus;
wire     [31:0] io_mp2_data_out_2_pinmux_mscbus;
wire     [31:0] io_mp2_dir_out_mscbus;
wire     [31:0] io_mp2_ds0_out_mscbus;
wire     [31:0] io_mp2_ds1_out_mscbus;
wire     [31:0] io_mp2_glitch_filter_bypass_out_mscbus;
wire     [63:0] io_mp2_glitch_filter_debounce_clk_sel_out_mscbus;
wire     [31:0] io_mp2_gpio_out_2_buf_mscbus;
wire     [31:0] io_mp2_gpio_out_en_2_buf_mscbus;
wire   [1023:0] io_mp2_in_function_en_out_mscbus;
wire     [31:0] io_mp2_in_termination_en_out_mscbus;
wire     [31:0] io_mp2_inena_out_mscbus;
wire     [31:0] io_mp2_lvds_en_ctrl_out_mscbus;
wire     [31:0] io_mp2_mode0_out_mscbus;
wire     [31:0] io_mp2_mode1_out_mscbus;
wire    [255:0] io_mp2_pes_en_out_mscbus;
wire     [31:0] io_mp2_pes_in_en_out_mscbus;
wire     [63:0] io_mp2_pes_safeval_out_mscbus;
wire    [159:0] io_mp2_pinmux_muxsel_out_mscbus;
wire     [31:0] io_mp2_pinmuxdata_2_gpio_mscbus;
wire     [31:0] io_mp2_pinmuxen_2_gpio_mscbus;
wire     [31:0] io_mp2_pull_en_out_mscbus;
wire     [31:0] io_mp2_pull_type_out_mscbus;
wire     [31:0] io_mp2_schmitt_out_mscbus;
wire     [31:0] io_mp2_slew_out_mscbus;
wire            io_reset_n;
wire     [31:0] io_vbusp_slv_address;
wire      [3:0] io_vbusp_slv_byten;
wire            io_vbusp_slv_dir;
wire      [1:0] io_vbusp_slv_dtype;
wire            io_vbusp_slv_emudbg;
wire      [1:0] io_vbusp_slv_priv;
wire      [7:0] io_vbusp_slv_privid;
wire     [31:0] io_vbusp_slv_rdatap;
wire            io_vbusp_slv_req;
wire     [11:0] io_vbusp_slv_routeid;
wire            io_vbusp_slv_rready;
wire      [2:0] io_vbusp_slv_rstatus;
wire            io_vbusp_slv_secure;
wire     [31:0] io_vbusp_slv_wdata;
wire            io_vbusp_slv_wready;
wire      [2:0] io_vbusp_slv_xcnt;
wire     [11:0] io_vbusp_slv_xid;
wire            jtag_tck;
wire            jtag_tdi;
wire            jtag_tdo;
wire            jtag_tdo_oe_n;
wire            jtag_tms;
wire            jtag_trst_n;
wire            o_porsn_frompad_reset_n;
wire            o_porsn_frompmm_pm_a_reset_n;
wire            o_porsn_frompmm_pm_b_reset_n;
wire            o_porsn_frompmm_pm_d_reset_n;
wire            o_porsn_pm_b_reset_n;
wire            o_porsn_sw_pm_a_reset_n;
wire            o_porsn_sw_pm_b_reset_n;
wire            o_porsn_sw_pm_d_reset_n;
wire            o_porsn_sw_streched_pm_a_reset_n;
wire            o_porsn_sw_streched_pm_b_reset_n;
wire            o_xrsn_frompad_reset_n;
wire            o_xrsn_pm_b_reset_n;
wire            o_xrsn_sw_fast_reset_n;
wire            o_xrsn_sw_streched_reset_n;
wire            pinmux_clock;
wire            pinmux_reset_n;
wire            sys_reset_n;
wire            xbar_clk_clock;
wire            xbar_rst_reset_n;

assign AP0_0_IO = AP0_IO;

assign AP0_1_IO = AP1_IO;

assign AP0_2_IO = AP2_IO;

assign AP0_3_IO = AP3_IO;

assign AP0_4_IO = AP4_IO;

assign AP0_5_IO = AP5_IO;

assign AP0_6_IO = AP6_IO;

assign AP0_7_IO = AP7_IO;

assign AP0_8_IO = AP8_IO;

assign AP0_9_IO = AP9_IO;

assign AP0_10_IO = AP10_IO;

assign AP0_11_IO = AP11_IO;

assign AP0_12_IO = AP12_IO;

assign AP0_13_IO = AP13_IO;

assign AP0_14_IO = AP14_IO;

assign AP0_15_IO = AP15_IO;

assign AP0_16_IO = AP16_IO;

assign AP0_17_IO = AP17_IO;

assign AP0_18_IO = AP18_IO;

assign AP0_19_IO = AP19_IO;

assign AP0_20_IO = AP20_IO;

assign AP0_21_IO = AP21_IO;

assign AP0_22_IO = AP22_IO;

assign AP0_23_IO = AP23_IO;

assign AP0_24_IO = AP24_IO;

assign AP0_25_IO = AP25_IO;

assign AP0_26_IO = AP26_IO;

assign AP0_27_IO = AP27_IO;

assign AP0_28_IO = AP28_IO;

assign AP0_29_IO = AP29_IO;

assign AP0_30_IO = AP30_IO;

assign AP0_31_IO = AP31_IO;

assign AP1_0_IO = AP32_IO;

assign AP1_1_IO = AP33_IO;

assign AP1_2_IO = AP34_IO;

assign AP1_3_IO = AP35_IO;

assign AP1_4_IO = AP36_IO;

assign AP1_5_IO = AP37_IO;

assign AP1_6_IO = AP38_IO;

assign AP1_7_IO = AP39_IO;

assign AP1_8_IO = AP40_IO;

assign AP1_9_IO = AP41_IO;

assign AP1_10_IO = AP42_IO;

assign AP1_11_IO = AP43_IO;

assign AP1_12_IO = AP44_IO;

assign AP1_13_IO = AP45_IO;

assign AP1_14_IO = AP46_IO;

assign AP1_15_IO = AP47_IO;

//-- Rev History
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
//-- Rev History
// documentation params
//  signal creation params
//  attribute params
//  determine the default value based on the polarity
assign jtag_tck = TCK_IO;

assign jtag_tms = TMS_IO;

assign jtag_tdi = TDI_IO;

assign TDO_IO = jtag_tdo;

assign o_xrsn_pm_b_reset_n = PWR_ON_RSTn_IO;

assign o_xrsn_sw_fast_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_frompmm_pm_d_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_pm_b_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_sw_pm_a_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_sw_pm_b_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_sw_pm_d_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_frompad_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_frompmm_pm_a_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_sw_streched_pm_a_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_frompmm_pm_b_reset_n = PWR_ON_RSTn_IO;

assign o_porsn_sw_streched_pm_b_reset_n = PWR_ON_RSTn_IO;

assign o_xrsn_frompad_reset_n = PWR_ON_RSTn_IO;

assign o_xrsn_sw_streched_reset_n = PWR_ON_RSTn_IO;

pinmux_wrapper I_b_pinmux_wrapper(
  .pinmux_clock(pinmux_clock),
  .pinmux_reset_n(pinmux_reset_n),
  .dp0_async_in_from_pad_mscbus(io_dp0_async_in_from_pad_mscbus),
  .dp0_gpio_out_2_buf_mscbus(io_dp0_gpio_out_2_buf_mscbus),
  .dp0_gpio_out_en_2_buf_mscbus(io_dp0_gpio_out_en_2_buf_mscbus),
  .dp0_pinmuxdata_2_gpio_mscbus(io_dp0_pinmuxdata_2_gpio_mscbus),
  .dp0_pinmuxen_2_gpio_mscbus(io_dp0_pinmuxen_2_gpio_mscbus),
  .dp0_data_out_2_pinmux_mscbus(io_dp0_data_out_2_pinmux_mscbus),
  .dp0_GP_DATA_IN_out_mscbus(io_dp0_GP_DATA_IN_out_mscbus),
  .dp0_pinmux_muxsel_out_mscbus(io_dp0_pinmux_muxsel_out_mscbus),
  .dp0_in_function_en_out_mscbus(io_dp0_in_function_en_out_mscbus),
  .dp0_amsel_out_mscbus(io_dp0_amsel_out_mscbus),
  .dp0_ds0_out_mscbus(io_dp0_ds0_out_mscbus),
  .dp0_ds1_out_mscbus(io_dp0_ds1_out_mscbus),
  .dp0_mode0_out_mscbus(io_dp0_mode0_out_mscbus),
  .dp0_mode1_out_mscbus(io_dp0_mode1_out_mscbus),
  .dp0_schmitt_out_mscbus(io_dp0_schmitt_out_mscbus),
  .dp0_slew_out_mscbus(io_dp0_slew_out_mscbus),
  .dp0_dir_out_mscbus(io_dp0_dir_out_mscbus),
  .dp0_pull_en_out_mscbus(io_dp0_pull_en_out_mscbus),
  .dp0_pull_type_out_mscbus(io_dp0_pull_type_out_mscbus),
  .dp0_glitch_filter_bypass_out_mscbus(io_dp0_glitch_filter_bypass_out_mscbus),
  .dp0_glitch_filter_debounce_clk_sel_out_mscbus(io_dp0_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp0_inena_out_mscbus(io_dp0_inena_out_mscbus),
  .dp0_pes_safeval_out_mscbus(io_dp0_pes_safeval_out_mscbus),
  .dp0_pes_in_en_out_mscbus(io_dp0_pes_in_en_out_mscbus),
  .dp0_pes_en_out_mscbus(io_dp0_pes_en_out_mscbus),
  .dp0_in_termination_en_out_mscbus(io_dp0_in_termination_en_out_mscbus),
  .dp0_lvds_en_ctrl_out_mscbus(io_dp0_lvds_en_ctrl_out_mscbus),
  .dp1_async_in_from_pad_mscbus(io_dp1_async_in_from_pad_mscbus),
  .dp1_gpio_out_2_buf_mscbus(io_dp1_gpio_out_2_buf_mscbus),
  .dp1_gpio_out_en_2_buf_mscbus(io_dp1_gpio_out_en_2_buf_mscbus),
  .dp1_pinmuxdata_2_gpio_mscbus(io_dp1_pinmuxdata_2_gpio_mscbus),
  .dp1_pinmuxen_2_gpio_mscbus(io_dp1_pinmuxen_2_gpio_mscbus),
  .dp1_data_out_2_pinmux_mscbus(io_dp1_data_out_2_pinmux_mscbus),
  .dp1_GP_DATA_IN_out_mscbus(io_dp1_GP_DATA_IN_out_mscbus),
  .dp1_pinmux_muxsel_out_mscbus(io_dp1_pinmux_muxsel_out_mscbus),
  .dp1_in_function_en_out_mscbus(io_dp1_in_function_en_out_mscbus),
  .dp1_amsel_out_mscbus(io_dp1_amsel_out_mscbus),
  .dp1_ds0_out_mscbus(io_dp1_ds0_out_mscbus),
  .dp1_ds1_out_mscbus(io_dp1_ds1_out_mscbus),
  .dp1_mode0_out_mscbus(io_dp1_mode0_out_mscbus),
  .dp1_mode1_out_mscbus(io_dp1_mode1_out_mscbus),
  .dp1_schmitt_out_mscbus(io_dp1_schmitt_out_mscbus),
  .dp1_slew_out_mscbus(io_dp1_slew_out_mscbus),
  .dp1_dir_out_mscbus(io_dp1_dir_out_mscbus),
  .dp1_pull_en_out_mscbus(io_dp1_pull_en_out_mscbus),
  .dp1_pull_type_out_mscbus(io_dp1_pull_type_out_mscbus),
  .dp1_glitch_filter_bypass_out_mscbus(io_dp1_glitch_filter_bypass_out_mscbus),
  .dp1_glitch_filter_debounce_clk_sel_out_mscbus(io_dp1_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp1_inena_out_mscbus(io_dp1_inena_out_mscbus),
  .dp1_pes_safeval_out_mscbus(io_dp1_pes_safeval_out_mscbus),
  .dp1_pes_in_en_out_mscbus(io_dp1_pes_in_en_out_mscbus),
  .dp1_pes_en_out_mscbus(io_dp1_pes_en_out_mscbus),
  .dp1_in_termination_en_out_mscbus(io_dp1_in_termination_en_out_mscbus),
  .dp1_lvds_en_ctrl_out_mscbus(io_dp1_lvds_en_ctrl_out_mscbus),
  .dp2_async_in_from_pad_mscbus(io_dp2_async_in_from_pad_mscbus),
  .dp2_gpio_out_2_buf_mscbus(io_dp2_gpio_out_2_buf_mscbus),
  .dp2_gpio_out_en_2_buf_mscbus(io_dp2_gpio_out_en_2_buf_mscbus),
  .dp2_pinmuxdata_2_gpio_mscbus(io_dp2_pinmuxdata_2_gpio_mscbus),
  .dp2_pinmuxen_2_gpio_mscbus(io_dp2_pinmuxen_2_gpio_mscbus),
  .dp2_data_out_2_pinmux_mscbus(io_dp2_data_out_2_pinmux_mscbus),
  .dp2_GP_DATA_IN_out_mscbus(io_dp2_GP_DATA_IN_out_mscbus),
  .dp2_pinmux_muxsel_out_mscbus(io_dp2_pinmux_muxsel_out_mscbus),
  .dp2_in_function_en_out_mscbus(io_dp2_in_function_en_out_mscbus),
  .dp2_amsel_out_mscbus(io_dp2_amsel_out_mscbus),
  .dp2_ds0_out_mscbus(io_dp2_ds0_out_mscbus),
  .dp2_ds1_out_mscbus(io_dp2_ds1_out_mscbus),
  .dp2_mode0_out_mscbus(io_dp2_mode0_out_mscbus),
  .dp2_mode1_out_mscbus(io_dp2_mode1_out_mscbus),
  .dp2_schmitt_out_mscbus(io_dp2_schmitt_out_mscbus),
  .dp2_slew_out_mscbus(io_dp2_slew_out_mscbus),
  .dp2_dir_out_mscbus(io_dp2_dir_out_mscbus),
  .dp2_pull_en_out_mscbus(io_dp2_pull_en_out_mscbus),
  .dp2_pull_type_out_mscbus(io_dp2_pull_type_out_mscbus),
  .dp2_glitch_filter_bypass_out_mscbus(io_dp2_glitch_filter_bypass_out_mscbus),
  .dp2_glitch_filter_debounce_clk_sel_out_mscbus(io_dp2_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp2_inena_out_mscbus(io_dp2_inena_out_mscbus),
  .dp2_pes_safeval_out_mscbus(io_dp2_pes_safeval_out_mscbus),
  .dp2_pes_in_en_out_mscbus(io_dp2_pes_in_en_out_mscbus),
  .dp2_pes_en_out_mscbus(io_dp2_pes_en_out_mscbus),
  .dp2_in_termination_en_out_mscbus(io_dp2_in_termination_en_out_mscbus),
  .dp2_lvds_en_ctrl_out_mscbus(io_dp2_lvds_en_ctrl_out_mscbus),
  .dp3_async_in_from_pad_mscbus(io_dp3_async_in_from_pad_mscbus),
  .dp3_gpio_out_2_buf_mscbus(io_dp3_gpio_out_2_buf_mscbus),
  .dp3_gpio_out_en_2_buf_mscbus(io_dp3_gpio_out_en_2_buf_mscbus),
  .dp3_pinmuxdata_2_gpio_mscbus(io_dp3_pinmuxdata_2_gpio_mscbus),
  .dp3_pinmuxen_2_gpio_mscbus(io_dp3_pinmuxen_2_gpio_mscbus),
  .dp3_data_out_2_pinmux_mscbus(io_dp3_data_out_2_pinmux_mscbus),
  .dp3_GP_DATA_IN_out_mscbus(io_dp3_GP_DATA_IN_out_mscbus),
  .dp3_pinmux_muxsel_out_mscbus(io_dp3_pinmux_muxsel_out_mscbus),
  .dp3_in_function_en_out_mscbus(io_dp3_in_function_en_out_mscbus),
  .dp3_amsel_out_mscbus(io_dp3_amsel_out_mscbus),
  .dp3_ds0_out_mscbus(io_dp3_ds0_out_mscbus),
  .dp3_ds1_out_mscbus(io_dp3_ds1_out_mscbus),
  .dp3_mode0_out_mscbus(io_dp3_mode0_out_mscbus),
  .dp3_mode1_out_mscbus(io_dp3_mode1_out_mscbus),
  .dp3_schmitt_out_mscbus(io_dp3_schmitt_out_mscbus),
  .dp3_slew_out_mscbus(io_dp3_slew_out_mscbus),
  .dp3_dir_out_mscbus(io_dp3_dir_out_mscbus),
  .dp3_pull_en_out_mscbus(io_dp3_pull_en_out_mscbus),
  .dp3_pull_type_out_mscbus(io_dp3_pull_type_out_mscbus),
  .dp3_glitch_filter_bypass_out_mscbus(io_dp3_glitch_filter_bypass_out_mscbus),
  .dp3_glitch_filter_debounce_clk_sel_out_mscbus(io_dp3_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp3_inena_out_mscbus(io_dp3_inena_out_mscbus),
  .dp3_pes_safeval_out_mscbus(io_dp3_pes_safeval_out_mscbus),
  .dp3_pes_in_en_out_mscbus(io_dp3_pes_in_en_out_mscbus),
  .dp3_pes_en_out_mscbus(io_dp3_pes_en_out_mscbus),
  .dp3_in_termination_en_out_mscbus(io_dp3_in_termination_en_out_mscbus),
  .dp3_lvds_en_ctrl_out_mscbus(io_dp3_lvds_en_ctrl_out_mscbus),
  .dp4_async_in_from_pad_mscbus(io_dp4_async_in_from_pad_mscbus),
  .dp4_gpio_out_2_buf_mscbus(io_dp4_gpio_out_2_buf_mscbus),
  .dp4_gpio_out_en_2_buf_mscbus(io_dp4_gpio_out_en_2_buf_mscbus),
  .dp4_pinmuxdata_2_gpio_mscbus(io_dp4_pinmuxdata_2_gpio_mscbus),
  .dp4_pinmuxen_2_gpio_mscbus(io_dp4_pinmuxen_2_gpio_mscbus),
  .dp4_data_out_2_pinmux_mscbus(io_dp4_data_out_2_pinmux_mscbus),
  .dp4_GP_DATA_IN_out_mscbus(io_dp4_GP_DATA_IN_out_mscbus),
  .dp4_pinmux_muxsel_out_mscbus(io_dp4_pinmux_muxsel_out_mscbus),
  .dp4_in_function_en_out_mscbus(io_dp4_in_function_en_out_mscbus),
  .dp4_amsel_out_mscbus(io_dp4_amsel_out_mscbus),
  .dp4_ds0_out_mscbus(io_dp4_ds0_out_mscbus),
  .dp4_ds1_out_mscbus(io_dp4_ds1_out_mscbus),
  .dp4_mode0_out_mscbus(io_dp4_mode0_out_mscbus),
  .dp4_mode1_out_mscbus(io_dp4_mode1_out_mscbus),
  .dp4_schmitt_out_mscbus(io_dp4_schmitt_out_mscbus),
  .dp4_slew_out_mscbus(io_dp4_slew_out_mscbus),
  .dp4_dir_out_mscbus(io_dp4_dir_out_mscbus),
  .dp4_pull_en_out_mscbus(io_dp4_pull_en_out_mscbus),
  .dp4_pull_type_out_mscbus(io_dp4_pull_type_out_mscbus),
  .dp4_glitch_filter_bypass_out_mscbus(io_dp4_glitch_filter_bypass_out_mscbus),
  .dp4_glitch_filter_debounce_clk_sel_out_mscbus(io_dp4_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp4_inena_out_mscbus(io_dp4_inena_out_mscbus),
  .dp4_pes_safeval_out_mscbus(io_dp4_pes_safeval_out_mscbus),
  .dp4_pes_in_en_out_mscbus(io_dp4_pes_in_en_out_mscbus),
  .dp4_pes_en_out_mscbus(io_dp4_pes_en_out_mscbus),
  .dp4_in_termination_en_out_mscbus(io_dp4_in_termination_en_out_mscbus),
  .dp4_lvds_en_ctrl_out_mscbus(io_dp4_lvds_en_ctrl_out_mscbus),
  .dp5_async_in_from_pad_mscbus(io_dp5_async_in_from_pad_mscbus),
  .dp5_gpio_out_2_buf_mscbus(io_dp5_gpio_out_2_buf_mscbus),
  .dp5_gpio_out_en_2_buf_mscbus(io_dp5_gpio_out_en_2_buf_mscbus),
  .dp5_pinmuxdata_2_gpio_mscbus(io_dp5_pinmuxdata_2_gpio_mscbus),
  .dp5_pinmuxen_2_gpio_mscbus(io_dp5_pinmuxen_2_gpio_mscbus),
  .dp5_data_out_2_pinmux_mscbus(io_dp5_data_out_2_pinmux_mscbus),
  .dp5_GP_DATA_IN_out_mscbus(io_dp5_GP_DATA_IN_out_mscbus),
  .dp5_pinmux_muxsel_out_mscbus(io_dp5_pinmux_muxsel_out_mscbus),
  .dp5_in_function_en_out_mscbus(io_dp5_in_function_en_out_mscbus),
  .dp5_amsel_out_mscbus(io_dp5_amsel_out_mscbus),
  .dp5_ds0_out_mscbus(io_dp5_ds0_out_mscbus),
  .dp5_ds1_out_mscbus(io_dp5_ds1_out_mscbus),
  .dp5_mode0_out_mscbus(io_dp5_mode0_out_mscbus),
  .dp5_mode1_out_mscbus(io_dp5_mode1_out_mscbus),
  .dp5_schmitt_out_mscbus(io_dp5_schmitt_out_mscbus),
  .dp5_slew_out_mscbus(io_dp5_slew_out_mscbus),
  .dp5_dir_out_mscbus(io_dp5_dir_out_mscbus),
  .dp5_pull_en_out_mscbus(io_dp5_pull_en_out_mscbus),
  .dp5_pull_type_out_mscbus(io_dp5_pull_type_out_mscbus),
  .dp5_glitch_filter_bypass_out_mscbus(io_dp5_glitch_filter_bypass_out_mscbus),
  .dp5_glitch_filter_debounce_clk_sel_out_mscbus(io_dp5_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp5_inena_out_mscbus(io_dp5_inena_out_mscbus),
  .dp5_pes_safeval_out_mscbus(io_dp5_pes_safeval_out_mscbus),
  .dp5_pes_in_en_out_mscbus(io_dp5_pes_in_en_out_mscbus),
  .dp5_pes_en_out_mscbus(io_dp5_pes_en_out_mscbus),
  .dp5_in_termination_en_out_mscbus(io_dp5_in_termination_en_out_mscbus),
  .dp5_lvds_en_ctrl_out_mscbus(io_dp5_lvds_en_ctrl_out_mscbus),
  .dp6_async_in_from_pad_mscbus(io_dp6_async_in_from_pad_mscbus),
  .dp6_gpio_out_2_buf_mscbus(io_dp6_gpio_out_2_buf_mscbus),
  .dp6_gpio_out_en_2_buf_mscbus(io_dp6_gpio_out_en_2_buf_mscbus),
  .dp6_pinmuxdata_2_gpio_mscbus(io_dp6_pinmuxdata_2_gpio_mscbus),
  .dp6_pinmuxen_2_gpio_mscbus(io_dp6_pinmuxen_2_gpio_mscbus),
  .dp6_data_out_2_pinmux_mscbus(io_dp6_data_out_2_pinmux_mscbus),
  .dp6_GP_DATA_IN_out_mscbus(io_dp6_GP_DATA_IN_out_mscbus),
  .dp6_pinmux_muxsel_out_mscbus(io_dp6_pinmux_muxsel_out_mscbus),
  .dp6_in_function_en_out_mscbus(io_dp6_in_function_en_out_mscbus),
  .dp6_amsel_out_mscbus(io_dp6_amsel_out_mscbus),
  .dp6_ds0_out_mscbus(io_dp6_ds0_out_mscbus),
  .dp6_ds1_out_mscbus(io_dp6_ds1_out_mscbus),
  .dp6_mode0_out_mscbus(io_dp6_mode0_out_mscbus),
  .dp6_mode1_out_mscbus(io_dp6_mode1_out_mscbus),
  .dp6_schmitt_out_mscbus(io_dp6_schmitt_out_mscbus),
  .dp6_slew_out_mscbus(io_dp6_slew_out_mscbus),
  .dp6_dir_out_mscbus(io_dp6_dir_out_mscbus),
  .dp6_pull_en_out_mscbus(io_dp6_pull_en_out_mscbus),
  .dp6_pull_type_out_mscbus(io_dp6_pull_type_out_mscbus),
  .dp6_glitch_filter_bypass_out_mscbus(io_dp6_glitch_filter_bypass_out_mscbus),
  .dp6_glitch_filter_debounce_clk_sel_out_mscbus(io_dp6_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp6_inena_out_mscbus(io_dp6_inena_out_mscbus),
  .dp6_pes_safeval_out_mscbus(io_dp6_pes_safeval_out_mscbus),
  .dp6_pes_in_en_out_mscbus(io_dp6_pes_in_en_out_mscbus),
  .dp6_pes_en_out_mscbus(io_dp6_pes_en_out_mscbus),
  .dp6_in_termination_en_out_mscbus(io_dp6_in_termination_en_out_mscbus),
  .dp6_lvds_en_ctrl_out_mscbus(io_dp6_lvds_en_ctrl_out_mscbus),
  .dp7_async_in_from_pad_mscbus(io_dp7_async_in_from_pad_mscbus),
  .dp7_gpio_out_2_buf_mscbus(io_dp7_gpio_out_2_buf_mscbus),
  .dp7_gpio_out_en_2_buf_mscbus(io_dp7_gpio_out_en_2_buf_mscbus),
  .dp7_pinmuxdata_2_gpio_mscbus(io_dp7_pinmuxdata_2_gpio_mscbus),
  .dp7_pinmuxen_2_gpio_mscbus(io_dp7_pinmuxen_2_gpio_mscbus),
  .dp7_data_out_2_pinmux_mscbus(io_dp7_data_out_2_pinmux_mscbus),
  .dp7_GP_DATA_IN_out_mscbus(io_dp7_GP_DATA_IN_out_mscbus),
  .dp7_pinmux_muxsel_out_mscbus(io_dp7_pinmux_muxsel_out_mscbus),
  .dp7_in_function_en_out_mscbus(io_dp7_in_function_en_out_mscbus),
  .dp7_amsel_out_mscbus(io_dp7_amsel_out_mscbus),
  .dp7_ds0_out_mscbus(io_dp7_ds0_out_mscbus),
  .dp7_ds1_out_mscbus(io_dp7_ds1_out_mscbus),
  .dp7_mode0_out_mscbus(io_dp7_mode0_out_mscbus),
  .dp7_mode1_out_mscbus(io_dp7_mode1_out_mscbus),
  .dp7_schmitt_out_mscbus(io_dp7_schmitt_out_mscbus),
  .dp7_slew_out_mscbus(io_dp7_slew_out_mscbus),
  .dp7_dir_out_mscbus(io_dp7_dir_out_mscbus),
  .dp7_pull_en_out_mscbus(io_dp7_pull_en_out_mscbus),
  .dp7_pull_type_out_mscbus(io_dp7_pull_type_out_mscbus),
  .dp7_glitch_filter_bypass_out_mscbus(io_dp7_glitch_filter_bypass_out_mscbus),
  .dp7_glitch_filter_debounce_clk_sel_out_mscbus(io_dp7_glitch_filter_debounce_clk_sel_out_mscbus),
  .dp7_inena_out_mscbus(io_dp7_inena_out_mscbus),
  .dp7_pes_safeval_out_mscbus(io_dp7_pes_safeval_out_mscbus),
  .dp7_pes_in_en_out_mscbus(io_dp7_pes_in_en_out_mscbus),
  .dp7_pes_en_out_mscbus(io_dp7_pes_en_out_mscbus),
  .dp7_in_termination_en_out_mscbus(io_dp7_in_termination_en_out_mscbus),
  .dp7_lvds_en_ctrl_out_mscbus(io_dp7_lvds_en_ctrl_out_mscbus),
  .mp0_async_in_from_pad_mscbus(io_mp0_async_in_from_pad_mscbus),
  .mp0_gpio_out_2_buf_mscbus(io_mp0_gpio_out_2_buf_mscbus),
  .mp0_gpio_out_en_2_buf_mscbus(io_mp0_gpio_out_en_2_buf_mscbus),
  .mp0_pinmuxdata_2_gpio_mscbus(io_mp0_pinmuxdata_2_gpio_mscbus),
  .mp0_pinmuxen_2_gpio_mscbus(io_mp0_pinmuxen_2_gpio_mscbus),
  .mp0_data_out_2_pinmux_mscbus(io_mp0_data_out_2_pinmux_mscbus),
  .mp0_GP_DATA_IN_out_mscbus(io_mp0_GP_DATA_IN_out_mscbus),
  .mp0_pinmux_muxsel_out_mscbus(io_mp0_pinmux_muxsel_out_mscbus),
  .mp0_in_function_en_out_mscbus(io_mp0_in_function_en_out_mscbus),
  .mp0_amsel_out_mscbus(io_mp0_amsel_out_mscbus),
  .mp0_ds0_out_mscbus(io_mp0_ds0_out_mscbus),
  .mp0_ds1_out_mscbus(io_mp0_ds1_out_mscbus),
  .mp0_mode0_out_mscbus(io_mp0_mode0_out_mscbus),
  .mp0_mode1_out_mscbus(io_mp0_mode1_out_mscbus),
  .mp0_schmitt_out_mscbus(io_mp0_schmitt_out_mscbus),
  .mp0_slew_out_mscbus(io_mp0_slew_out_mscbus),
  .mp0_dir_out_mscbus(io_mp0_dir_out_mscbus),
  .mp0_pull_en_out_mscbus(io_mp0_pull_en_out_mscbus),
  .mp0_pull_type_out_mscbus(io_mp0_pull_type_out_mscbus),
  .mp0_glitch_filter_bypass_out_mscbus(io_mp0_glitch_filter_bypass_out_mscbus),
  .mp0_glitch_filter_debounce_clk_sel_out_mscbus(io_mp0_glitch_filter_debounce_clk_sel_out_mscbus),
  .mp0_inena_out_mscbus(io_mp0_inena_out_mscbus),
  .mp0_pes_safeval_out_mscbus(io_mp0_pes_safeval_out_mscbus),
  .mp0_pes_in_en_out_mscbus(io_mp0_pes_in_en_out_mscbus),
  .mp0_pes_en_out_mscbus(io_mp0_pes_en_out_mscbus),
  .mp0_in_termination_en_out_mscbus(io_mp0_in_termination_en_out_mscbus),
  .mp0_lvds_en_ctrl_out_mscbus(io_mp0_lvds_en_ctrl_out_mscbus),
  .mp1_async_in_from_pad_mscbus(io_mp1_async_in_from_pad_mscbus),
  .mp1_gpio_out_2_buf_mscbus(io_mp1_gpio_out_2_buf_mscbus),
  .mp1_gpio_out_en_2_buf_mscbus(io_mp1_gpio_out_en_2_buf_mscbus),
  .mp1_pinmuxdata_2_gpio_mscbus(io_mp1_pinmuxdata_2_gpio_mscbus),
  .mp1_pinmuxen_2_gpio_mscbus(io_mp1_pinmuxen_2_gpio_mscbus),
  .mp1_data_out_2_pinmux_mscbus(io_mp1_data_out_2_pinmux_mscbus),
  .mp1_GP_DATA_IN_out_mscbus(io_mp1_GP_DATA_IN_out_mscbus),
  .mp1_pinmux_muxsel_out_mscbus(io_mp1_pinmux_muxsel_out_mscbus),
  .mp1_in_function_en_out_mscbus(io_mp1_in_function_en_out_mscbus),
  .mp1_amsel_out_mscbus(io_mp1_amsel_out_mscbus),
  .mp1_ds0_out_mscbus(io_mp1_ds0_out_mscbus),
  .mp1_ds1_out_mscbus(io_mp1_ds1_out_mscbus),
  .mp1_mode0_out_mscbus(io_mp1_mode0_out_mscbus),
  .mp1_mode1_out_mscbus(io_mp1_mode1_out_mscbus),
  .mp1_schmitt_out_mscbus(io_mp1_schmitt_out_mscbus),
  .mp1_slew_out_mscbus(io_mp1_slew_out_mscbus),
  .mp1_dir_out_mscbus(io_mp1_dir_out_mscbus),
  .mp1_pull_en_out_mscbus(io_mp1_pull_en_out_mscbus),
  .mp1_pull_type_out_mscbus(io_mp1_pull_type_out_mscbus),
  .mp1_glitch_filter_bypass_out_mscbus(io_mp1_glitch_filter_bypass_out_mscbus),
  .mp1_glitch_filter_debounce_clk_sel_out_mscbus(io_mp1_glitch_filter_debounce_clk_sel_out_mscbus),
  .mp1_inena_out_mscbus(io_mp1_inena_out_mscbus),
  .mp1_pes_safeval_out_mscbus(io_mp1_pes_safeval_out_mscbus),
  .mp1_pes_in_en_out_mscbus(io_mp1_pes_in_en_out_mscbus),
  .mp1_pes_en_out_mscbus(io_mp1_pes_en_out_mscbus),
  .mp1_in_termination_en_out_mscbus(io_mp1_in_termination_en_out_mscbus),
  .mp1_lvds_en_ctrl_out_mscbus(io_mp1_lvds_en_ctrl_out_mscbus),
  .mp2_async_in_from_pad_mscbus(io_mp2_async_in_from_pad_mscbus),
  .mp2_gpio_out_2_buf_mscbus(io_mp2_gpio_out_2_buf_mscbus),
  .mp2_gpio_out_en_2_buf_mscbus(io_mp2_gpio_out_en_2_buf_mscbus),
  .mp2_pinmuxdata_2_gpio_mscbus(io_mp2_pinmuxdata_2_gpio_mscbus),
  .mp2_pinmuxen_2_gpio_mscbus(io_mp2_pinmuxen_2_gpio_mscbus),
  .mp2_data_out_2_pinmux_mscbus(io_mp2_data_out_2_pinmux_mscbus),
  .mp2_GP_DATA_IN_out_mscbus(io_mp2_GP_DATA_IN_out_mscbus),
  .mp2_pinmux_muxsel_out_mscbus(io_mp2_pinmux_muxsel_out_mscbus),
  .mp2_in_function_en_out_mscbus(io_mp2_in_function_en_out_mscbus),
  .mp2_amsel_out_mscbus(io_mp2_amsel_out_mscbus),
  .mp2_ds0_out_mscbus(io_mp2_ds0_out_mscbus),
  .mp2_ds1_out_mscbus(io_mp2_ds1_out_mscbus),
  .mp2_mode0_out_mscbus(io_mp2_mode0_out_mscbus),
  .mp2_mode1_out_mscbus(io_mp2_mode1_out_mscbus),
  .mp2_schmitt_out_mscbus(io_mp2_schmitt_out_mscbus),
  .mp2_slew_out_mscbus(io_mp2_slew_out_mscbus),
  .mp2_dir_out_mscbus(io_mp2_dir_out_mscbus),
  .mp2_pull_en_out_mscbus(io_mp2_pull_en_out_mscbus),
  .mp2_pull_type_out_mscbus(io_mp2_pull_type_out_mscbus),
  .mp2_glitch_filter_bypass_out_mscbus(io_mp2_glitch_filter_bypass_out_mscbus),
  .mp2_glitch_filter_debounce_clk_sel_out_mscbus(io_mp2_glitch_filter_debounce_clk_sel_out_mscbus),
  .mp2_inena_out_mscbus(io_mp2_inena_out_mscbus),
  .mp2_pes_safeval_out_mscbus(io_mp2_pes_safeval_out_mscbus),
  .mp2_pes_in_en_out_mscbus(io_mp2_pes_in_en_out_mscbus),
  .mp2_pes_en_out_mscbus(io_mp2_pes_en_out_mscbus),
  .mp2_in_termination_en_out_mscbus(io_mp2_in_termination_en_out_mscbus),
  .mp2_lvds_en_ctrl_out_mscbus(io_mp2_lvds_en_ctrl_out_mscbus),
  .ap0_async_in_from_pad_mscbus(io_ap0_async_in_from_pad_mscbus),
  .ap0_gpio_out_2_buf_mscbus(io_ap0_gpio_out_2_buf_mscbus),
  .ap0_gpio_out_en_2_buf_mscbus(io_ap0_gpio_out_en_2_buf_mscbus),
  .ap0_pinmuxdata_2_gpio_mscbus(io_ap0_pinmuxdata_2_gpio_mscbus),
  .ap0_pinmuxen_2_gpio_mscbus(io_ap0_pinmuxen_2_gpio_mscbus),
  .ap0_data_out_2_pinmux_mscbus(io_ap0_data_out_2_pinmux_mscbus),
  .ap0_GP_DATA_IN_out_mscbus(io_ap0_GP_DATA_IN_out_mscbus),
  .ap0_pinmux_muxsel_out_mscbus(io_ap0_pinmux_muxsel_out_mscbus),
  .ap0_in_function_en_out_mscbus(io_ap0_in_function_en_out_mscbus),
  .ap0_amsel_out_mscbus(io_ap0_amsel_out_mscbus),
  .ap0_ds0_out_mscbus(io_ap0_ds0_out_mscbus),
  .ap0_ds1_out_mscbus(io_ap0_ds1_out_mscbus),
  .ap0_mode0_out_mscbus(io_ap0_mode0_out_mscbus),
  .ap0_mode1_out_mscbus(io_ap0_mode1_out_mscbus),
  .ap0_schmitt_out_mscbus(io_ap0_schmitt_out_mscbus),
  .ap0_slew_out_mscbus(io_ap0_slew_out_mscbus),
  .ap0_dir_out_mscbus(io_ap0_dir_out_mscbus),
  .ap0_pull_en_out_mscbus(io_ap0_pull_en_out_mscbus),
  .ap0_pull_type_out_mscbus(io_ap0_pull_type_out_mscbus),
  .ap0_glitch_filter_bypass_out_mscbus(io_ap0_glitch_filter_bypass_out_mscbus),
  .ap0_glitch_filter_debounce_clk_sel_out_mscbus(io_ap0_glitch_filter_debounce_clk_sel_out_mscbus),
  .ap0_inena_out_mscbus(io_ap0_inena_out_mscbus),
  .ap0_pes_safeval_out_mscbus(io_ap0_pes_safeval_out_mscbus),
  .ap0_pes_in_en_out_mscbus(io_ap0_pes_in_en_out_mscbus),
  .ap0_pes_en_out_mscbus(io_ap0_pes_en_out_mscbus),
  .ap0_in_termination_en_out_mscbus(io_ap0_in_termination_en_out_mscbus),
  .ap0_lvds_en_ctrl_out_mscbus(io_ap0_lvds_en_ctrl_out_mscbus),
  .ap1_async_in_from_pad_mscbus(io_ap1_async_in_from_pad_mscbus),
  .ap1_gpio_out_2_buf_mscbus(io_ap1_gpio_out_2_buf_mscbus),
  .ap1_gpio_out_en_2_buf_mscbus(io_ap1_gpio_out_en_2_buf_mscbus),
  .ap1_pinmuxdata_2_gpio_mscbus(io_ap1_pinmuxdata_2_gpio_mscbus),
  .ap1_pinmuxen_2_gpio_mscbus(io_ap1_pinmuxen_2_gpio_mscbus),
  .ap1_data_out_2_pinmux_mscbus(io_ap1_data_out_2_pinmux_mscbus),
  .ap1_GP_DATA_IN_out_mscbus(io_ap1_GP_DATA_IN_out_mscbus),
  .ap1_pinmux_muxsel_out_mscbus(io_ap1_pinmux_muxsel_out_mscbus),
  .ap1_in_function_en_out_mscbus(io_ap1_in_function_en_out_mscbus),
  .ap1_amsel_out_mscbus(io_ap1_amsel_out_mscbus),
  .ap1_ds0_out_mscbus(io_ap1_ds0_out_mscbus),
  .ap1_ds1_out_mscbus(io_ap1_ds1_out_mscbus),
  .ap1_mode0_out_mscbus(io_ap1_mode0_out_mscbus),
  .ap1_mode1_out_mscbus(io_ap1_mode1_out_mscbus),
  .ap1_schmitt_out_mscbus(io_ap1_schmitt_out_mscbus),
  .ap1_slew_out_mscbus(io_ap1_slew_out_mscbus),
  .ap1_dir_out_mscbus(io_ap1_dir_out_mscbus),
  .ap1_pull_en_out_mscbus(io_ap1_pull_en_out_mscbus),
  .ap1_pull_type_out_mscbus(io_ap1_pull_type_out_mscbus),
  .ap1_glitch_filter_bypass_out_mscbus(io_ap1_glitch_filter_bypass_out_mscbus),
  .ap1_glitch_filter_debounce_clk_sel_out_mscbus(io_ap1_glitch_filter_debounce_clk_sel_out_mscbus),
  .ap1_inena_out_mscbus(io_ap1_inena_out_mscbus),
  .ap1_pes_safeval_out_mscbus(io_ap1_pes_safeval_out_mscbus),
  .ap1_pes_in_en_out_mscbus(io_ap1_pes_in_en_out_mscbus),
  .ap1_pes_en_out_mscbus(io_ap1_pes_en_out_mscbus),
  .ap1_in_termination_en_out_mscbus(io_ap1_in_termination_en_out_mscbus),
  .ap1_lvds_en_ctrl_out_mscbus(io_ap1_lvds_en_ctrl_out_mscbus),
  .DP0_0_IO(DP0_0_IO),
  .DP0_1_IO(DP0_1_IO),
  .DP0_2_IO(DP0_2_IO),
  .DP0_3_IO(DP0_3_IO),
  .DP0_4_IO(DP0_4_IO),
  .DP0_5_IO(DP0_5_IO),
  .DP0_6_IO(DP0_6_IO),
  .DP0_7_IO(DP0_7_IO),
  .DP0_8_IO(DP0_8_IO),
  .DP0_9_IO(DP0_9_IO),
  .DP0_10_IO(DP0_10_IO),
  .DP0_11_IO(DP0_11_IO),
  .DP0_12_IO(DP0_12_IO),
  .DP0_13_IO(DP0_13_IO),
  .DP0_14_IO(DP0_14_IO),
  .DP0_15_IO(DP0_15_IO),
  .DP0_16_IO(DP0_16_IO),
  .DP0_17_IO(DP0_17_IO),
  .DP0_18_IO(DP0_18_IO),
  .DP0_19_IO(DP0_19_IO),
  .DP0_20_IO(DP0_20_IO),
  .DP0_21_IO(DP0_21_IO),
  .DP0_22_IO(DP0_22_IO),
  .DP0_23_IO(DP0_23_IO),
  .DP0_24_IO(DP0_24_IO),
  .DP0_25_IO(DP0_25_IO),
  .DP0_26_IO(DP0_26_IO),
  .DP0_27_IO(DP0_27_IO),
  .DP0_28_IO(DP0_28_IO),
  .DP0_29_IO(DP0_29_IO),
  .DP0_30_IO(DP0_30_IO),
  .DP0_31_IO(DP0_31_IO),
  .DP1_0_IO(DP1_0_IO),
  .DP1_1_IO(DP1_1_IO),
  .DP1_2_IO(DP1_2_IO),
  .DP1_3_IO(DP1_3_IO),
  .DP1_4_IO(DP1_4_IO),
  .DP1_5_IO(DP1_5_IO),
  .DP1_6_IO(DP1_6_IO),
  .DP1_7_IO(DP1_7_IO),
  .DP1_8_IO(DP1_8_IO),
  .DP1_9_IO(DP1_9_IO),
  .DP1_10_IO(DP1_10_IO),
  .DP1_11_IO(DP1_11_IO),
  .DP1_12_IO(DP1_12_IO),
  .DP1_13_IO(DP1_13_IO),
  .DP1_14_IO(DP1_14_IO),
  .DP1_15_IO(DP1_15_IO),
  .DP1_16_IO(DP1_16_IO),
  .DP1_17_IO(DP1_17_IO),
  .DP1_18_IO(DP1_18_IO),
  .DP1_19_IO(DP1_19_IO),
  .DP1_20_IO(DP1_20_IO),
  .DP1_21_IO(DP1_21_IO),
  .DP1_22_IO(DP1_22_IO),
  .DP1_23_IO(DP1_23_IO),
  .DP1_24_IO(DP1_24_IO),
  .DP1_25_IO(DP1_25_IO),
  .DP1_26_IO(DP1_26_IO),
  .DP1_27_IO(DP1_27_IO),
  .DP1_28_IO(DP1_28_IO),
  .DP1_29_IO(DP1_29_IO),
  .DP1_30_IO(DP1_30_IO),
  .DP1_31_IO(DP1_31_IO),
  .DP2_0_IO(DP2_0_IO),
  .DP2_1_IO(DP2_1_IO),
  .DP2_2_IO(DP2_2_IO),
  .DP2_3_IO(DP2_3_IO),
  .DP2_4_IO(DP2_4_IO),
  .DP2_5_IO(DP2_5_IO),
  .DP2_6_IO(DP2_6_IO),
  .DP2_7_IO(DP2_7_IO),
  .DP2_8_IO(DP2_8_IO),
  .DP2_9_IO(DP2_9_IO),
  .DP2_10_IO(DP2_10_IO),
  .DP2_11_IO(DP2_11_IO),
  .DP2_12_IO(DP2_12_IO),
  .DP2_13_IO(DP2_13_IO),
  .DP2_14_IO(DP2_14_IO),
  .DP2_15_IO(DP2_15_IO),
  .DP2_16_IO(DP2_16_IO),
  .DP2_17_IO(DP2_17_IO),
  .DP2_18_IO(DP2_18_IO),
  .DP2_19_IO(DP2_19_IO),
  .DP2_20_IO(DP2_20_IO),
  .DP2_21_IO(DP2_21_IO),
  .DP2_22_IO(DP2_22_IO),
  .DP2_23_IO(DP2_23_IO),
  .DP2_24_IO(DP2_24_IO),
  .DP2_25_IO(DP2_25_IO),
  .DP2_26_IO(DP2_26_IO),
  .DP2_27_IO(DP2_27_IO),
  .DP2_28_IO(DP2_28_IO),
  .DP2_29_IO(DP2_29_IO),
  .DP2_30_IO(DP2_30_IO),
  .DP2_31_IO(DP2_31_IO),
  .DP3_0_IO(DP3_0_IO),
  .DP3_1_IO(DP3_1_IO),
  .DP3_2_IO(DP3_2_IO),
  .DP3_3_IO(DP3_3_IO),
  .DP3_4_IO(DP3_4_IO),
  .DP3_5_IO(DP3_5_IO),
  .DP3_6_IO(DP3_6_IO),
  .DP3_7_IO(DP3_7_IO),
  .DP3_8_IO(DP3_8_IO),
  .DP3_9_IO(DP3_9_IO),
  .DP3_10_IO(DP3_10_IO),
  .DP3_11_IO(DP3_11_IO),
  .DP3_12_IO(DP3_12_IO),
  .DP3_13_IO(DP3_13_IO),
  .DP3_14_IO(DP3_14_IO),
  .DP3_15_IO(DP3_15_IO),
  .DP3_16_IO(DP3_16_IO),
  .DP3_17_IO(DP3_17_IO),
  .DP3_18_IO(DP3_18_IO),
  .DP3_19_IO(DP3_19_IO),
  .DP3_20_IO(DP3_20_IO),
  .DP3_21_IO(DP3_21_IO),
  .DP3_22_IO(DP3_22_IO),
  .DP3_23_IO(DP3_23_IO),
  .DP3_24_IO(DP3_24_IO),
  .DP3_25_IO(DP3_25_IO),
  .DP3_26_IO(DP3_26_IO),
  .DP3_27_IO(DP3_27_IO),
  .DP3_28_IO(DP3_28_IO),
  .DP3_29_IO(DP3_29_IO),
  .DP3_30_IO(DP3_30_IO),
  .DP3_31_IO(DP3_31_IO),
  .DP4_0_IO(DP4_0_IO),
  .DP4_1_IO(DP4_1_IO),
  .DP4_2_IO(DP4_2_IO),
  .DP4_3_IO(DP4_3_IO),
  .DP4_4_IO(DP4_4_IO),
  .DP4_5_IO(DP4_5_IO),
  .DP4_6_IO(DP4_6_IO),
  .DP4_7_IO(DP4_7_IO),
  .DP4_8_IO(DP4_8_IO),
  .DP4_9_IO(DP4_9_IO),
  .DP4_10_IO(DP4_10_IO),
  .DP4_11_IO(DP4_11_IO),
  .DP4_12_IO(DP4_12_IO),
  .DP4_13_IO(DP4_13_IO),
  .DP4_14_IO(DP4_14_IO),
  .DP4_15_IO(DP4_15_IO),
  .DP4_16_IO(DP4_16_IO),
  .DP4_17_IO(DP4_17_IO),
  .DP4_18_IO(DP4_18_IO),
  .DP4_19_IO(DP4_19_IO),
  .DP4_20_IO(DP4_20_IO),
  .DP4_21_IO(DP4_21_IO),
  .DP4_22_IO(DP4_22_IO),
  .DP4_23_IO(DP4_23_IO),
  .DP4_24_IO(DP4_24_IO),
  .DP4_25_IO(DP4_25_IO),
  .DP4_26_IO(DP4_26_IO),
  .DP4_27_IO(DP4_27_IO),
  .DP4_28_IO(DP4_28_IO),
  .DP4_29_IO(DP4_29_IO),
  .DP4_30_IO(DP4_30_IO),
  .DP4_31_IO(DP4_31_IO),
  .DP5_0_IO(DP5_0_IO),
  .DP5_1_IO(DP5_1_IO),
  .DP5_2_IO(DP5_2_IO),
  .DP5_3_IO(DP5_3_IO),
  .DP5_4_IO(DP5_4_IO),
  .DP5_5_IO(DP5_5_IO),
  .DP5_6_IO(DP5_6_IO),
  .DP5_7_IO(DP5_7_IO),
  .DP5_8_IO(DP5_8_IO),
  .DP5_9_IO(DP5_9_IO),
  .DP5_10_IO(DP5_10_IO),
  .DP5_11_IO(DP5_11_IO),
  .DP5_12_IO(DP5_12_IO),
  .DP5_13_IO(DP5_13_IO),
  .DP5_14_IO(DP5_14_IO),
  .DP5_15_IO(DP5_15_IO),
  .DP5_16_IO(DP5_16_IO),
  .DP5_17_IO(DP5_17_IO),
  .DP5_18_IO(DP5_18_IO),
  .DP5_19_IO(DP5_19_IO),
  .DP5_20_IO(DP5_20_IO),
  .DP5_21_IO(DP5_21_IO),
  .DP5_22_IO(DP5_22_IO),
  .DP5_23_IO(DP5_23_IO),
  .DP5_24_IO(DP5_24_IO),
  .DP5_25_IO(DP5_25_IO),
  .DP5_26_IO(DP5_26_IO),
  .DP5_27_IO(DP5_27_IO),
  .DP5_28_IO(DP5_28_IO),
  .DP5_29_IO(DP5_29_IO),
  .DP5_30_IO(DP5_30_IO),
  .DP5_31_IO(DP5_31_IO),
  .DP6_0_IO(DP6_0_IO),
  .DP6_1_IO(DP6_1_IO),
  .DP6_2_IO(DP6_2_IO),
  .DP6_3_IO(DP6_3_IO),
  .DP6_4_IO(DP6_4_IO),
  .DP6_5_IO(DP6_5_IO),
  .DP6_6_IO(DP6_6_IO),
  .DP6_7_IO(DP6_7_IO),
  .DP6_8_IO(DP6_8_IO),
  .DP6_9_IO(DP6_9_IO),
  .DP6_10_IO(DP6_10_IO),
  .DP6_11_IO(DP6_11_IO),
  .DP6_12_IO(DP6_12_IO),
  .DP6_13_IO(DP6_13_IO),
  .DP6_14_IO(DP6_14_IO),
  .DP6_15_IO(DP6_15_IO),
  .DP6_16_IO(DP6_16_IO),
  .DP6_17_IO(DP6_17_IO),
  .DP6_18_IO(DP6_18_IO),
  .DP6_19_IO(DP6_19_IO),
  .DP6_20_IO(DP6_20_IO),
  .DP6_21_IO(DP6_21_IO),
  .DP6_22_IO(DP6_22_IO),
  .DP6_23_IO(DP6_23_IO),
  .DP6_24_IO(DP6_24_IO),
  .DP6_25_IO(DP6_25_IO),
  .DP6_26_IO(DP6_26_IO),
  .DP6_27_IO(DP6_27_IO),
  .DP7_0_IO(DP7_0_IO),
  .DP7_1_IO(DP7_1_IO),
  .DP7_2_IO(DP7_2_IO),
  .DP7_3_IO(DP7_3_IO),
  .DP7_4_IO(DP7_4_IO),
  .DP7_5_IO(DP7_5_IO),
  .DP7_6_IO(DP7_6_IO),
  .DP7_7_IO(DP7_7_IO),
  .DP7_8_IO(DP7_8_IO),
  .DP7_9_IO(DP7_9_IO),
  .DP7_10_IO(DP7_10_IO),
  .DP7_11_IO(DP7_11_IO),
  .DP7_12_IO(DP7_12_IO),
  .DP7_13_IO(DP7_13_IO),
  .DP7_14_IO(DP7_14_IO),
  .DP7_15_IO(DP7_15_IO),
  .MP0_0_IO(MP0_0_IO),
  .MP0_1_IO(MP0_1_IO),
  .MP0_2_IO(MP0_2_IO),
  .MP0_3_IO(MP0_3_IO),
  .MP0_4_IO(MP0_4_IO),
  .MP0_5_IO(MP0_5_IO),
  .MP0_6_IO(MP0_6_IO),
  .MP0_7_IO(MP0_7_IO),
  .MP0_8_IO(MP0_8_IO),
  .MP0_9_IO(MP0_9_IO),
  .MP0_10_IO(MP0_10_IO),
  .MP0_11_IO(MP0_11_IO),
  .MP0_12_IO(MP0_12_IO),
  .MP0_13_IO(MP0_13_IO),
  .MP0_14_IO(MP0_14_IO),
  .MP0_15_IO(MP0_15_IO),
  .MP0_16_IO(MP0_16_IO),
  .MP0_17_IO(MP0_17_IO),
  .MP0_18_IO(MP0_18_IO),
  .MP0_19_IO(MP0_19_IO),
  .MP0_20_IO(MP0_20_IO),
  .MP0_21_IO(MP0_21_IO),
  .MP0_22_IO(MP0_22_IO),
  .MP0_23_IO(MP0_23_IO),
  .MP0_24_IO(MP0_24_IO),
  .MP0_25_IO(MP0_25_IO),
  .MP0_26_IO(MP0_26_IO),
  .MP0_27_IO(MP0_27_IO),
  .MP0_28_IO(MP0_28_IO),
  .MP0_29_IO(MP0_29_IO),
  .MP0_30_IO(MP0_30_IO),
  .MP0_31_IO(MP0_31_IO),
  .MP1_0_IO(MP1_0_IO),
  .MP1_1_IO(MP1_1_IO),
  .MP1_2_IO(MP1_2_IO),
  .MP1_3_IO(MP1_3_IO),
  .MP1_4_IO(MP1_4_IO),
  .MP1_5_IO(MP1_5_IO),
  .MP1_6_IO(MP1_6_IO),
  .MP1_7_IO(MP1_7_IO),
  .MP1_8_IO(MP1_8_IO),
  .MP1_9_IO(MP1_9_IO),
  .MP1_10_IO(MP1_10_IO),
  .MP1_11_IO(MP1_11_IO),
  .MP1_12_IO(MP1_12_IO),
  .MP1_13_IO(MP1_13_IO),
  .MP1_14_IO(MP1_14_IO),
  .MP1_15_IO(MP1_15_IO),
  .MP2_0_IO(MP2_0_IO),
  .MP2_1_IO(MP2_1_IO),
  .MP2_2_IO(MP2_2_IO),
  .MP2_3_IO(MP2_3_IO),
  .MP2_4_IO(MP2_4_IO),
  .MP2_5_IO(MP2_5_IO),
  .MP2_6_IO(MP2_6_IO),
  .MP2_7_IO(MP2_7_IO),
  .MP2_8_IO(MP2_8_IO),
  .MP2_9_IO(MP2_9_IO),
  .MP2_10_IO(MP2_10_IO),
  .MP2_11_IO(MP2_11_IO),
  .MP2_12_IO(MP2_12_IO),
  .MP2_13_IO(MP2_13_IO),
  .MP2_14_IO(MP2_14_IO),
  .MP2_15_IO(MP2_15_IO),
  .AP0_0_IO(AP0_0_IO),
  .AP0_1_IO(AP0_1_IO),
  .AP0_2_IO(AP0_2_IO),
  .AP0_3_IO(AP0_3_IO),
  .AP0_4_IO(AP0_4_IO),
  .AP0_5_IO(AP0_5_IO),
  .AP0_6_IO(AP0_6_IO),
  .AP0_7_IO(AP0_7_IO),
  .AP0_8_IO(AP0_8_IO),
  .AP0_9_IO(AP0_9_IO),
  .AP0_10_IO(AP0_10_IO),
  .AP0_11_IO(AP0_11_IO),
  .AP0_12_IO(AP0_12_IO),
  .AP0_13_IO(AP0_13_IO),
  .AP0_14_IO(AP0_14_IO),
  .AP0_15_IO(AP0_15_IO),
  .AP0_16_IO(AP0_16_IO),
  .AP0_17_IO(AP0_17_IO),
  .AP0_18_IO(AP0_18_IO),
  .AP0_19_IO(AP0_19_IO),
  .AP0_20_IO(AP0_20_IO),
  .AP0_21_IO(AP0_21_IO),
  .AP0_22_IO(AP0_22_IO),
  .AP0_23_IO(AP0_23_IO),
  .AP0_24_IO(AP0_24_IO),
  .AP0_25_IO(AP0_25_IO),
  .AP0_26_IO(AP0_26_IO),
  .AP0_27_IO(AP0_27_IO),
  .AP0_28_IO(AP0_28_IO),
  .AP0_29_IO(AP0_29_IO),
  .AP0_30_IO(AP0_30_IO),
  .AP0_31_IO(AP0_31_IO),
  .AP1_0_IO(AP1_0_IO),
  .AP1_1_IO(AP1_1_IO),
  .AP1_2_IO(AP1_2_IO),
  .AP1_3_IO(AP1_3_IO),
  .AP1_4_IO(AP1_4_IO),
  .AP1_5_IO(AP1_5_IO),
  .AP1_6_IO(AP1_6_IO),
  .AP1_7_IO(AP1_7_IO),
  .AP1_8_IO(AP1_8_IO),
  .AP1_9_IO(AP1_9_IO),
  .AP1_10_IO(AP1_10_IO),
  .AP1_11_IO(AP1_11_IO),
  .AP1_12_IO(AP1_12_IO),
  .AP1_13_IO(AP1_13_IO),
  .AP1_14_IO(AP1_14_IO),
  .AP1_15_IO(AP1_15_IO)
);

// RTL Assignments for DP ports
// Auto-generated - Do not edit
// Assignments for DP0_0
assign DP0_0_in_mux_peripheral_mscbus[1] = io_CAN0_txd;

assign DP0_0_in_mux_en_mscbus[1] = 1'b0;

assign DP0_0_in_mux_peripheral_mscbus[3] = io_EPWM0_a_o;

assign DP0_0_in_mux_en_mscbus[3] = io_EPWM0_a_oen;

assign DP0_0_in_mux_peripheral_mscbus[4] = io_SPI8PICO_out;

assign DP0_0_in_mux_en_mscbus[4] = io_SPI8PICO_oen;

assign DP0_0_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR6_intr;

assign DP0_0_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP0_0
// Assignments for DP0_1
assign DP0_1_in_mux_peripheral_mscbus[2] = io_EPWM0_b_o;

assign DP0_1_in_mux_en_mscbus[2] = io_EPWM0_b_oen;

assign DP0_1_in_mux_peripheral_mscbus[3] = io_OUTPUTXBAR7_intr;

assign DP0_1_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP0_1
assign io_CAN0_rxd = DP0_1_out_demux_peripheral_mscbus[1];

assign io_SPI8POCI_in = DP0_1_out_demux_peripheral_mscbus[2];

// Assignments for DP0_10
assign DP0_10_in_mux_peripheral_mscbus[1] = io_FSI0TX_ck;

assign DP0_10_in_mux_en_mscbus[1] = 1'b0;

assign DP0_10_in_mux_peripheral_mscbus[3] = io_EPWM5_a_o;

assign DP0_10_in_mux_en_mscbus[3] = io_EPWM5_a_oen;

assign DP0_10_in_mux_peripheral_mscbus[4] = io_SPI9CS1_out;

assign DP0_10_in_mux_en_mscbus[4] = io_SPI9CS1_oen;

// Assignments for DP0_10
// Assignments for DP0_11
assign DP0_11_in_mux_peripheral_mscbus[1] = io_FSI0TX_d0;

assign DP0_11_in_mux_en_mscbus[1] = 1'b0;

assign DP0_11_in_mux_peripheral_mscbus[3] = io_EPWM5_b_o;

assign DP0_11_in_mux_en_mscbus[3] = io_EPWM5_b_oen;

assign DP0_11_in_mux_peripheral_mscbus[4] = io_SPI9CS2_out;

assign DP0_11_in_mux_en_mscbus[4] = io_SPI9CS2_oen;

// Assignments for DP0_11
// Assignments for DP0_12
assign DP0_12_in_mux_peripheral_mscbus[1] = io_FSI0TX_d1;

assign DP0_12_in_mux_en_mscbus[1] = 1'b0;

assign DP0_12_in_mux_peripheral_mscbus[3] = io_EPWM6_a_o;

assign DP0_12_in_mux_en_mscbus[3] = io_EPWM6_a_oen;

assign DP0_12_in_mux_peripheral_mscbus[4] = io_SPI9CS3_out;

assign DP0_12_in_mux_en_mscbus[4] = io_SPI9CS3_oen;

// Assignments for DP0_12
// Assignments for DP0_13
assign DP0_13_in_mux_peripheral_mscbus[2] = io_EPWM6_b_o;

assign DP0_13_in_mux_en_mscbus[2] = io_EPWM6_b_oen;

assign DP0_13_in_mux_peripheral_mscbus[3] = io_FSI0TX_ck;

assign DP0_13_in_mux_en_mscbus[3] = 1'b0;

assign DP0_13_in_mux_peripheral_mscbus[5] = io_SPI9CS4_out;

assign DP0_13_in_mux_en_mscbus[5] = io_SPI9CS4_oen;

// Assignments for DP0_13
assign io_FSI0RX_ck = DP0_13_out_demux_peripheral_mscbus[1];

// Assignments for DP0_14
assign DP0_14_in_mux_peripheral_mscbus[2] = io_EPWM7_a_o;

assign DP0_14_in_mux_en_mscbus[2] = io_EPWM7_a_oen;

assign DP0_14_in_mux_peripheral_mscbus[3] = io_FSI0TX_d0;

assign DP0_14_in_mux_en_mscbus[3] = 1'b0;

assign DP0_14_in_mux_peripheral_mscbus[5] = io_SPI2CLK_clock;

assign DP0_14_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP0_14
assign io_FSI0RX_d0 = DP0_14_out_demux_peripheral_mscbus[1];

// Assignments for DP0_15
assign DP0_15_in_mux_peripheral_mscbus[2] = io_EPWM7_b_o;

assign DP0_15_in_mux_en_mscbus[2] = io_EPWM7_b_oen;

assign DP0_15_in_mux_peripheral_mscbus[3] = io_FSI0TX_d1;

assign DP0_15_in_mux_en_mscbus[3] = 1'b0;

assign DP0_15_in_mux_peripheral_mscbus[5] = io_SPI2PICO_out;

assign DP0_15_in_mux_en_mscbus[5] = io_SPI2PICO_oen;

// Assignments for DP0_15
assign io_FSI0RX_d1 = DP0_15_out_demux_peripheral_mscbus[1];

// Assignments for DP0_16
assign DP0_16_in_mux_peripheral_mscbus[3] = io_EPWM8_a_o;

assign DP0_16_in_mux_en_mscbus[3] = io_EPWM8_a_oen;

// Assignments for DP0_16
assign io_FSI0RX_ck = DP0_16_out_demux_peripheral_mscbus[2];

assign io_SPI2POCI_in = DP0_16_out_demux_peripheral_mscbus[3];

// Assignments for DP0_17
assign DP0_17_in_mux_peripheral_mscbus[3] = io_EPWM8_b_o;

assign DP0_17_in_mux_en_mscbus[3] = io_EPWM8_b_oen;

assign DP0_17_in_mux_peripheral_mscbus[5] = io_SPI2CS0_out;

assign DP0_17_in_mux_en_mscbus[5] = io_SPI2CS0_oen;

// Assignments for DP0_17
assign io_FSI0RX_d0 = DP0_17_out_demux_peripheral_mscbus[2];

// Assignments for DP0_18
assign DP0_18_in_mux_peripheral_mscbus[3] = io_EPWM9_a_o;

assign DP0_18_in_mux_en_mscbus[3] = io_EPWM9_a_oen;

assign DP0_18_in_mux_peripheral_mscbus[5] = io_SPI2CS1_out;

assign DP0_18_in_mux_en_mscbus[5] = io_SPI2CS1_oen;

// Assignments for DP0_18
assign io_FSI0RX_d1 = DP0_18_out_demux_peripheral_mscbus[2];

// Assignments for DP0_19
assign DP0_19_in_mux_peripheral_mscbus[3] = io_EPWM9_b_o;

assign DP0_19_in_mux_en_mscbus[3] = io_EPWM9_b_oen;

assign DP0_19_in_mux_peripheral_mscbus[4] = io_FSI1TX_ck;

assign DP0_19_in_mux_en_mscbus[4] = 1'b0;

assign DP0_19_in_mux_peripheral_mscbus[6] = io_SPI2CS2_out;

assign DP0_19_in_mux_en_mscbus[6] = io_SPI2CS2_oen;

// Assignments for DP0_19
// Assignments for DP0_2
assign DP0_2_in_mux_peripheral_mscbus[1] = io_CAN1_txd;

assign DP0_2_in_mux_en_mscbus[1] = 1'b0;

assign DP0_2_in_mux_peripheral_mscbus[3] = io_EPWM1_a_o;

assign DP0_2_in_mux_en_mscbus[3] = io_EPWM1_a_oen;

assign DP0_2_in_mux_peripheral_mscbus[4] = io_SPI8CS0_out;

assign DP0_2_in_mux_en_mscbus[4] = io_SPI8CS0_oen;

assign DP0_2_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR8_intr;

assign DP0_2_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP0_2
// Assignments for DP0_20
assign DP0_20_in_mux_peripheral_mscbus[1] = io_LIN0_txd;

assign DP0_20_in_mux_en_mscbus[1] = io_LIN0_tr_en;

assign DP0_20_in_mux_peripheral_mscbus[3] = io_EPWM10_a_o;

assign DP0_20_in_mux_en_mscbus[3] = io_EPWM10_b_oen;

assign DP0_20_in_mux_peripheral_mscbus[4] = io_FSI1TX_d0;

assign DP0_20_in_mux_en_mscbus[4] = 1'b0;

assign DP0_20_in_mux_peripheral_mscbus[6] = io_SPI2CS3_out;

assign DP0_20_in_mux_en_mscbus[6] = io_SPI2CS3_oen;

// Assignments for DP0_20
// Assignments for DP0_21
assign DP0_21_in_mux_peripheral_mscbus[2] = io_EPWM10_b_o;

assign DP0_21_in_mux_en_mscbus[2] = io_EPWM10_b_oen;

assign DP0_21_in_mux_peripheral_mscbus[3] = io_FSI1TX_d1;

assign DP0_21_in_mux_en_mscbus[3] = 1'b0;

assign DP0_21_in_mux_peripheral_mscbus[5] = io_LIN4_txd;

assign DP0_21_in_mux_en_mscbus[5] = io_LIN4_tr_en;

// Assignments for DP0_21
assign io_LIN0_rxd = DP0_21_out_demux_peripheral_mscbus[1];

// Assignments for DP0_22
assign DP0_22_in_mux_peripheral_mscbus[1] = io_LIN1_txd;

assign DP0_22_in_mux_en_mscbus[1] = io_LIN1_tr_en;

assign DP0_22_in_mux_peripheral_mscbus[3] = io_EPWM11_a_o;

assign DP0_22_in_mux_en_mscbus[3] = io_EPWM11_a_oen;

// Assignments for DP0_22
assign io_FSI1RX_ck = DP0_22_out_demux_peripheral_mscbus[1];

assign io_LIN4_rxd = DP0_22_out_demux_peripheral_mscbus[2];

// Assignments for DP0_23
assign DP0_23_in_mux_peripheral_mscbus[1] = io_SPI7CS3_out;

assign DP0_23_in_mux_en_mscbus[1] = io_SPI7CS3_oen;

assign DP0_23_in_mux_peripheral_mscbus[2] = io_EPWM11_b_o;

assign DP0_23_in_mux_en_mscbus[2] = io_EPWM11_b_oen;

assign DP0_23_in_mux_peripheral_mscbus[4] = io_LIN5_txd;

assign DP0_23_in_mux_en_mscbus[4] = io_LIN5_tr_en;

// Assignments for DP0_23
assign io_LIN1_rxd = DP0_23_out_demux_peripheral_mscbus[1];

assign io_FSI1RX_d0 = DP0_23_out_demux_peripheral_mscbus[2];

// Assignments for DP0_24
assign DP0_24_in_mux_peripheral_mscbus[1] = io_LIN2_txd;

assign DP0_24_in_mux_en_mscbus[1] = io_LIN2_tr_en;

assign DP0_24_in_mux_peripheral_mscbus[2] = io_SPI7CLK_clock;

assign DP0_24_in_mux_en_mscbus[2] = 1'b0;

assign DP0_24_in_mux_peripheral_mscbus[3] = io_EPWM12_a_o;

assign DP0_24_in_mux_en_mscbus[3] = io_EPWM12_a_oen;

// Assignments for DP0_24
assign io_FSI1RX_d1 = DP0_24_out_demux_peripheral_mscbus[1];

assign io_LIN5_rxd = DP0_24_out_demux_peripheral_mscbus[2];

// Assignments for DP0_25
assign DP0_25_in_mux_peripheral_mscbus[1] = io_SPI7PICO_out;

assign DP0_25_in_mux_en_mscbus[1] = io_SPI7PICO_oen;

assign DP0_25_in_mux_peripheral_mscbus[2] = io_EPWM12_b_o;

assign DP0_25_in_mux_en_mscbus[2] = io_EPWM12_b_oen;

assign DP0_25_in_mux_peripheral_mscbus[3] = io_FSI2TX_ck;

assign DP0_25_in_mux_en_mscbus[3] = 1'b0;

assign DP0_25_in_mux_peripheral_mscbus[5] = io_SPI5CS4_out;

assign DP0_25_in_mux_en_mscbus[5] = io_SPI5CS4_oen;

// Assignments for DP0_25
assign io_LIN2_rxd = DP0_25_out_demux_peripheral_mscbus[1];

// Assignments for DP0_26
assign DP0_26_in_mux_peripheral_mscbus[1] = io_LIN3_txd;

assign DP0_26_in_mux_en_mscbus[1] = io_LIN3_tr_en;

assign DP0_26_in_mux_peripheral_mscbus[2] = io_EPWM13_a_o;

assign DP0_26_in_mux_en_mscbus[2] = io_EPWM13_a_oen;

assign DP0_26_in_mux_peripheral_mscbus[3] = io_FSI2TX_d0;

assign DP0_26_in_mux_en_mscbus[3] = 1'b0;

assign DP0_26_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR0_intr;

assign DP0_26_in_mux_en_mscbus[4] = 1'b0;

assign DP0_26_in_mux_peripheral_mscbus[5] = io_SPI5CS5_out;

assign DP0_26_in_mux_en_mscbus[5] = io_SPI5CS5_oen;

// Assignments for DP0_26
assign io_SPI7POCI_in = DP0_26_out_demux_peripheral_mscbus[1];

// Assignments for DP0_27
assign DP0_27_in_mux_peripheral_mscbus[1] = io_SPI7CS0_out;

assign DP0_27_in_mux_en_mscbus[1] = io_SPI7CS0_oen;

assign DP0_27_in_mux_peripheral_mscbus[2] = io_EPWM13_b_o;

assign DP0_27_in_mux_en_mscbus[2] = io_EPWM13_b_oen;

assign DP0_27_in_mux_peripheral_mscbus[3] = io_FSI2TX_d1;

assign DP0_27_in_mux_en_mscbus[3] = 1'b0;

assign DP0_27_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR1_intr;

assign DP0_27_in_mux_en_mscbus[4] = 1'b0;

assign DP0_27_in_mux_peripheral_mscbus[5] = io_SPI9CS5_out;

assign DP0_27_in_mux_en_mscbus[5] = io_SPI9CS5_oen;

// Assignments for DP0_27
assign io_LIN3_rxd = DP0_27_out_demux_peripheral_mscbus[1];

// Assignments for DP0_28
assign DP0_28_in_mux_peripheral_mscbus[1] = io_UART0_tx;

assign DP0_28_in_mux_en_mscbus[1] = 1'b0;

assign DP0_28_in_mux_peripheral_mscbus[2] = io_SPI7CS1_out;

assign DP0_28_in_mux_en_mscbus[2] = io_SPI7CS1_oen;

assign DP0_28_in_mux_peripheral_mscbus[3] = io_EPWM14_a_o;

assign DP0_28_in_mux_en_mscbus[3] = io_EPWM14_a_oen;

assign DP0_28_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR2_intr;

assign DP0_28_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_28
assign io_FSI2RX_ck = DP0_28_out_demux_peripheral_mscbus[1];

// Assignments for DP0_29
assign DP0_29_in_mux_peripheral_mscbus[1] = io_SPI7CS2_out;

assign DP0_29_in_mux_en_mscbus[1] = io_SPI7CS2_oen;

assign DP0_29_in_mux_peripheral_mscbus[2] = io_EPWM14_b_o;

assign DP0_29_in_mux_en_mscbus[2] = io_EPWM14_b_oen;

assign DP0_29_in_mux_peripheral_mscbus[3] = io_OUTPUTXBAR3_intr;

assign DP0_29_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP0_29
assign io_UART0_rx = DP0_29_out_demux_peripheral_mscbus[1];

assign io_FSI2RX_d0 = DP0_29_out_demux_peripheral_mscbus[2];

// Assignments for DP0_3
assign DP0_3_in_mux_peripheral_mscbus[2] = io_EPWM1_b_o;

assign DP0_3_in_mux_en_mscbus[2] = io_EPWM1_a_oen;

assign DP0_3_in_mux_peripheral_mscbus[3] = io_SPI8CS1_out;

assign DP0_3_in_mux_en_mscbus[3] = io_SPI8CS1_oen;

assign DP0_3_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR9_intr;

assign DP0_3_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_3
assign io_CAN1_rxd = DP0_3_out_demux_peripheral_mscbus[1];

// Assignments for DP0_30
assign DP0_30_in_mux_peripheral_mscbus[1] = io_SPI5CLK_clock;

assign DP0_30_in_mux_en_mscbus[1] = 1'b0;

assign DP0_30_in_mux_peripheral_mscbus[2] = io_EPWM15_a_o;

assign DP0_30_in_mux_en_mscbus[2] = io_EPWM15_a_oen;

assign DP0_30_in_mux_peripheral_mscbus[3] = io_OUTPUTXBAR4_intr;

assign DP0_30_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP0_30
assign io_SENT0_rxd_i = DP0_30_out_demux_peripheral_mscbus[1];

assign io_FSI2RX_d1 = DP0_30_out_demux_peripheral_mscbus[2];

// Assignments for DP0_31
assign DP0_31_in_mux_peripheral_mscbus[1] = io_SPI5PICO_out;

assign DP0_31_in_mux_en_mscbus[1] = io_SPI5PICO_oen;

assign DP0_31_in_mux_peripheral_mscbus[2] = io_EPWM15_b_o;

assign DP0_31_in_mux_en_mscbus[2] = io_EPWM15_b_oen;

assign DP0_31_in_mux_peripheral_mscbus[3] = io_FSI3TX_ck;

assign DP0_31_in_mux_en_mscbus[3] = 1'b0;

assign DP0_31_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR5_intr;

assign DP0_31_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_31
assign io_SENT1_rxd_i = DP0_31_out_demux_peripheral_mscbus[1];

// Assignments for DP0_4
assign DP0_4_in_mux_peripheral_mscbus[1] = io_CAN2_txd;

assign DP0_4_in_mux_en_mscbus[1] = 1'b0;

assign DP0_4_in_mux_peripheral_mscbus[3] = io_EPWM2_a_o;

assign DP0_4_in_mux_en_mscbus[3] = io_EPWM2_a_oen;

assign DP0_4_in_mux_peripheral_mscbus[4] = io_SPI8CS2_out;

assign DP0_4_in_mux_en_mscbus[4] = io_SPI8CS2_oen;

assign DP0_4_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR10_intr;

assign DP0_4_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP0_4
// Assignments for DP0_5
assign DP0_5_in_mux_peripheral_mscbus[2] = io_EPWM2_b_o;

assign DP0_5_in_mux_en_mscbus[2] = io_EPWM2_b_oen;

assign DP0_5_in_mux_peripheral_mscbus[3] = io_SPI8CS3_out;

assign DP0_5_in_mux_en_mscbus[3] = io_SPI8CS3_oen;

assign DP0_5_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR11_intr;

assign DP0_5_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_5
assign io_CAN2_rxd = DP0_5_out_demux_peripheral_mscbus[1];

// Assignments for DP0_6
assign DP0_6_in_mux_peripheral_mscbus[1] = io_CAN3_txd;

assign DP0_6_in_mux_en_mscbus[1] = 1'b0;

assign DP0_6_in_mux_peripheral_mscbus[3] = io_EPWM3_a_o;

assign DP0_6_in_mux_en_mscbus[3] = io_EPWM3_a_oen;

assign DP0_6_in_mux_peripheral_mscbus[4] = io_SPI9CLK_clock;

assign DP0_6_in_mux_en_mscbus[4] = 1'b0;

assign DP0_6_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR12_intr;

assign DP0_6_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP0_6
// Assignments for DP0_7
assign DP0_7_in_mux_peripheral_mscbus[2] = io_EPWM3_b_o;

assign DP0_7_in_mux_en_mscbus[2] = io_EPWM3_b_oen;

assign DP0_7_in_mux_peripheral_mscbus[3] = io_SPI9PICO_out;

assign DP0_7_in_mux_en_mscbus[3] = io_SPI9PICO_oen;

assign DP0_7_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR13_intr;

assign DP0_7_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_7
assign io_CAN3_rxd = DP0_7_out_demux_peripheral_mscbus[1];

// Assignments for DP0_8
assign DP0_8_in_mux_peripheral_mscbus[1] = io_CAN4_txd;

assign DP0_8_in_mux_en_mscbus[1] = 1'b0;

assign DP0_8_in_mux_peripheral_mscbus[3] = io_EPWM4_a_o;

assign DP0_8_in_mux_en_mscbus[3] = io_EPWM4_a_oen;

assign DP0_8_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR14_intr;

assign DP0_8_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_8
assign io_SPI9POCI_in = DP0_8_out_demux_peripheral_mscbus[1];

// Assignments for DP0_9
assign DP0_9_in_mux_peripheral_mscbus[2] = io_EPWM4_b_o;

assign DP0_9_in_mux_en_mscbus[2] = io_EPWM4_b_oen;

assign DP0_9_in_mux_peripheral_mscbus[3] = io_SPI9CS0_out;

assign DP0_9_in_mux_en_mscbus[3] = io_SPI9CS0_oen;

assign DP0_9_in_mux_peripheral_mscbus[4] = io_OUTPUTXBAR15_intr;

assign DP0_9_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP0_9
assign io_CAN4_rxd = DP0_9_out_demux_peripheral_mscbus[1];

// Assignments for DP1_0
assign DP1_0_in_mux_peripheral_mscbus[1] = io_EPWM0_a_o;

assign DP1_0_in_mux_en_mscbus[1] = io_EPWM0_a_oen;

assign DP1_0_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR0_intr;

assign DP1_0_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_0
assign io_SDFM0_i_clock1 = DP1_0_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_ck = DP1_0_out_demux_peripheral_mscbus[2];

// Assignments for DP1_1
assign DP1_1_in_mux_peripheral_mscbus[1] = io_EPWM0_b_o;

assign DP1_1_in_mux_en_mscbus[1] = io_EPWM0_b_oen;

assign DP1_1_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR1_intr;

assign DP1_1_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_1
assign io_SDFM0_i_datain1 = DP1_1_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_d0 = DP1_1_out_demux_peripheral_mscbus[2];

// Assignments for DP1_10
assign DP1_10_in_mux_peripheral_mscbus[1] = io_EPWM5_a_o;

assign DP1_10_in_mux_en_mscbus[1] = io_EPWM5_a_oen;

assign DP1_10_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR10_intr;

assign DP1_10_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_10
assign io_SDFM5_i_clock1 = DP1_10_out_demux_peripheral_mscbus[1];

// Assignments for DP1_11
assign DP1_11_in_mux_peripheral_mscbus[1] = io_EPWM5_b_o;

assign DP1_11_in_mux_en_mscbus[1] = io_EPWM5_b_oen;

assign DP1_11_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR11_intr;

assign DP1_11_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_11
assign io_SDFM5_i_datain1 = DP1_11_out_demux_peripheral_mscbus[1];

// Assignments for DP1_12
assign DP1_12_in_mux_peripheral_mscbus[1] = io_EPWM6_a_o;

assign DP1_12_in_mux_en_mscbus[1] = io_EPWM6_a_oen;

assign DP1_12_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR12_intr;

assign DP1_12_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_12
assign io_SDFM6_i_clock1 = DP1_12_out_demux_peripheral_mscbus[1];

// Assignments for DP1_13
assign DP1_13_in_mux_peripheral_mscbus[1] = io_EPWM6_b_o;

assign DP1_13_in_mux_en_mscbus[1] = io_EPWM6_b_oen;

assign DP1_13_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR13_intr;

assign DP1_13_in_mux_en_mscbus[2] = 1'b0;

assign DP1_13_in_mux_peripheral_mscbus[3] = io_UART0_tx;

assign DP1_13_in_mux_en_mscbus[3] = 1'b0;

assign DP1_13_in_mux_peripheral_mscbus[4] = io_LIN0_txd;

assign DP1_13_in_mux_en_mscbus[4] = io_LIN0_tr_en;

// Assignments for DP1_13
assign io_SDFM6_i_datain1 = DP1_13_out_demux_peripheral_mscbus[1];

// Assignments for DP1_14
assign DP1_14_in_mux_peripheral_mscbus[1] = io_EPWM7_a_o;

assign DP1_14_in_mux_en_mscbus[1] = io_EPWM7_a_oen;

assign DP1_14_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR14_intr;

assign DP1_14_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_14
assign io_SDFM7_i_clock1 = DP1_14_out_demux_peripheral_mscbus[1];

assign io_UART0_rx = DP1_14_out_demux_peripheral_mscbus[2];

assign io_LIN0_rxd = DP1_14_out_demux_peripheral_mscbus[3];

// Assignments for DP1_15
assign DP1_15_in_mux_peripheral_mscbus[1] = io_EPWM7_b_o;

assign DP1_15_in_mux_en_mscbus[1] = io_EPWM7_b_oen;

assign DP1_15_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR15_intr;

assign DP1_15_in_mux_en_mscbus[2] = 1'b0;

assign DP1_15_in_mux_peripheral_mscbus[3] = io_SPI8CLK_clock;

assign DP1_15_in_mux_en_mscbus[3] = 1'b0;

assign DP1_15_in_mux_peripheral_mscbus[4] = io_LIN1_txd;

assign DP1_15_in_mux_en_mscbus[4] = io_LIN1_tr_en;

// Assignments for DP1_15
assign io_SDFM7_i_datain1 = DP1_15_out_demux_peripheral_mscbus[1];

// Assignments for DP1_16
assign DP1_16_in_mux_peripheral_mscbus[1] = io_EPWM8_a_o;

assign DP1_16_in_mux_en_mscbus[1] = io_EPWM8_a_oen;

assign DP1_16_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR0_intr;

assign DP1_16_in_mux_en_mscbus[2] = 1'b0;

assign DP1_16_in_mux_peripheral_mscbus[3] = io_SPI8PICO_out;

assign DP1_16_in_mux_en_mscbus[3] = io_SPI8PICO_oen;

// Assignments for DP1_16
assign io_SDFM8_i_clock1 = DP1_16_out_demux_peripheral_mscbus[1];

assign io_LIN1_rxd = DP1_16_out_demux_peripheral_mscbus[2];

// Assignments for DP1_17
assign DP1_17_in_mux_peripheral_mscbus[1] = io_EPWM8_b_o;

assign DP1_17_in_mux_en_mscbus[1] = io_EPWM8_b_oen;

assign DP1_17_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR1_intr;

assign DP1_17_in_mux_en_mscbus[2] = 1'b0;

assign DP1_17_in_mux_peripheral_mscbus[3] = io_LIN2_txd;

assign DP1_17_in_mux_en_mscbus[3] = io_LIN2_tr_en;

// Assignments for DP1_17
assign io_SDFM8_i_datain1 = DP1_17_out_demux_peripheral_mscbus[1];

assign io_SPI8POCI_in = DP1_17_out_demux_peripheral_mscbus[2];

// Assignments for DP1_18
assign DP1_18_in_mux_peripheral_mscbus[1] = io_EPWM9_a_o;

assign DP1_18_in_mux_en_mscbus[1] = io_EPWM9_a_oen;

assign DP1_18_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR2_intr;

assign DP1_18_in_mux_en_mscbus[2] = 1'b0;

assign DP1_18_in_mux_peripheral_mscbus[3] = io_SPI8CS0_out;

assign DP1_18_in_mux_en_mscbus[3] = io_SPI8CS0_oen;

// Assignments for DP1_18
assign io_SDFM9_i_clock1 = DP1_18_out_demux_peripheral_mscbus[1];

assign io_LIN2_rxd = DP1_18_out_demux_peripheral_mscbus[2];

// Assignments for DP1_19
assign DP1_19_in_mux_peripheral_mscbus[1] = io_EPWM9_b_o;

assign DP1_19_in_mux_en_mscbus[1] = io_EPWM9_b_oen;

assign DP1_19_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR3_intr;

assign DP1_19_in_mux_en_mscbus[2] = 1'b0;

assign DP1_19_in_mux_peripheral_mscbus[3] = io_SPI8CS1_out;

assign DP1_19_in_mux_en_mscbus[3] = io_SPI8CS1_oen;

assign DP1_19_in_mux_peripheral_mscbus[4] = io_LIN3_txd;

assign DP1_19_in_mux_en_mscbus[4] = io_LIN3_tr_en;

// Assignments for DP1_19
assign io_SDFM9_i_datain1 = DP1_19_out_demux_peripheral_mscbus[1];

// Assignments for DP1_2
assign DP1_2_in_mux_peripheral_mscbus[1] = io_EPWM1_a_o;

assign DP1_2_in_mux_en_mscbus[1] = io_EPWM1_a_oen;

assign DP1_2_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR2_intr;

assign DP1_2_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_2
assign io_SDFM1_i_clock1 = DP1_2_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_d1 = DP1_2_out_demux_peripheral_mscbus[2];

// Assignments for DP1_20
assign DP1_20_in_mux_peripheral_mscbus[1] = io_EPWM10_a_o;

assign DP1_20_in_mux_en_mscbus[1] = io_EPWM10_b_oen;

assign DP1_20_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR4_intr;

assign DP1_20_in_mux_en_mscbus[2] = 1'b0;

assign DP1_20_in_mux_peripheral_mscbus[3] = io_SPI8CS2_out;

assign DP1_20_in_mux_en_mscbus[3] = io_SPI8CS2_oen;

// Assignments for DP1_20
assign io_SDFM10_i_clock1 = DP1_20_out_demux_peripheral_mscbus[1];

assign io_LIN3_rxd = DP1_20_out_demux_peripheral_mscbus[2];

// Assignments for DP1_21
assign DP1_21_in_mux_peripheral_mscbus[1] = io_EPWM10_b_o;

assign DP1_21_in_mux_en_mscbus[1] = io_EPWM10_b_oen;

assign DP1_21_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR5_intr;

assign DP1_21_in_mux_en_mscbus[2] = 1'b0;

assign DP1_21_in_mux_peripheral_mscbus[3] = io_SPI8CS3_out;

assign DP1_21_in_mux_en_mscbus[3] = io_SPI8CS3_oen;

assign DP1_21_in_mux_peripheral_mscbus[4] = io_SPI4CS4_out;

assign DP1_21_in_mux_en_mscbus[4] = io_SPI4CS4_oen;

// Assignments for DP1_21
assign io_SDFM10_i_datain1 = DP1_21_out_demux_peripheral_mscbus[1];

// Assignments for DP1_22
assign DP1_22_in_mux_peripheral_mscbus[1] = io_EPWM11_a_o;

assign DP1_22_in_mux_en_mscbus[1] = io_EPWM11_a_oen;

assign DP1_22_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR6_intr;

assign DP1_22_in_mux_en_mscbus[2] = 1'b0;

assign DP1_22_in_mux_peripheral_mscbus[3] = io_SPI2CLK_clock;

assign DP1_22_in_mux_en_mscbus[3] = 1'b0;

assign DP1_22_in_mux_peripheral_mscbus[4] = io_SPI4CS5_out;

assign DP1_22_in_mux_en_mscbus[4] = io_SPI4CS5_oen;

// Assignments for DP1_22
assign io_SDFM11_i_clock1 = DP1_22_out_demux_peripheral_mscbus[1];

// Assignments for DP1_23
assign DP1_23_in_mux_peripheral_mscbus[1] = io_EPWM11_b_o;

assign DP1_23_in_mux_en_mscbus[1] = io_EPWM11_b_oen;

assign DP1_23_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR7_intr;

assign DP1_23_in_mux_en_mscbus[2] = 1'b0;

assign DP1_23_in_mux_peripheral_mscbus[3] = io_SPI2PICO_out;

assign DP1_23_in_mux_en_mscbus[3] = io_SPI2PICO_oen;

// Assignments for DP1_23
assign io_SDFM11_i_datain1 = DP1_23_out_demux_peripheral_mscbus[1];

// Assignments for DP1_24
assign DP1_24_in_mux_peripheral_mscbus[1] = io_EPWM12_a_o;

assign DP1_24_in_mux_en_mscbus[1] = io_EPWM12_a_oen;

assign DP1_24_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR8_intr;

assign DP1_24_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_24
assign io_SPI2POCI_in = DP1_24_out_demux_peripheral_mscbus[1];

// Assignments for DP1_25
assign DP1_25_in_mux_peripheral_mscbus[1] = io_EPWM12_b_o;

assign DP1_25_in_mux_en_mscbus[1] = io_EPWM12_b_oen;

assign DP1_25_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR9_intr;

assign DP1_25_in_mux_en_mscbus[2] = 1'b0;

assign DP1_25_in_mux_peripheral_mscbus[4] = io_SPI2CS0_out;

assign DP1_25_in_mux_en_mscbus[4] = io_SPI2CS0_oen;

// Assignments for DP1_25
// Assignments for DP1_26
assign DP1_26_in_mux_peripheral_mscbus[1] = io_EPWM13_a_o;

assign DP1_26_in_mux_en_mscbus[1] = io_EPWM13_a_oen;

assign DP1_26_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR10_intr;

assign DP1_26_in_mux_en_mscbus[2] = 1'b0;

assign DP1_26_in_mux_peripheral_mscbus[4] = io_SPI2CS1_out;

assign DP1_26_in_mux_en_mscbus[4] = io_SPI2CS1_oen;

// Assignments for DP1_26
// Assignments for DP1_27
assign DP1_27_in_mux_peripheral_mscbus[1] = io_EPWM13_b_o;

assign DP1_27_in_mux_en_mscbus[1] = io_EPWM13_b_oen;

assign DP1_27_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR11_intr;

assign DP1_27_in_mux_en_mscbus[2] = 1'b0;

assign DP1_27_in_mux_peripheral_mscbus[4] = io_SPI2CS2_out;

assign DP1_27_in_mux_en_mscbus[4] = io_SPI2CS2_oen;

// Assignments for DP1_27
// Assignments for DP1_28
assign DP1_28_in_mux_peripheral_mscbus[1] = io_EPWM14_a_o;

assign DP1_28_in_mux_en_mscbus[1] = io_EPWM14_a_oen;

assign DP1_28_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR12_intr;

assign DP1_28_in_mux_en_mscbus[2] = 1'b0;

assign DP1_28_in_mux_peripheral_mscbus[4] = io_SPI2CS3_out;

assign DP1_28_in_mux_en_mscbus[4] = io_SPI2CS3_oen;

// Assignments for DP1_28
// Assignments for DP1_29
assign DP1_29_in_mux_peripheral_mscbus[1] = io_EPWM14_b_o;

assign DP1_29_in_mux_en_mscbus[1] = io_EPWM14_b_oen;

assign DP1_29_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR13_intr;

assign DP1_29_in_mux_en_mscbus[2] = 1'b0;

assign DP1_29_in_mux_peripheral_mscbus[4] = io_SPI3CLK_clock;

assign DP1_29_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP1_29
// Assignments for DP1_3
assign DP1_3_in_mux_peripheral_mscbus[1] = io_EPWM1_b_o;

assign DP1_3_in_mux_en_mscbus[1] = io_EPWM1_a_oen;

assign DP1_3_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR3_intr;

assign DP1_3_in_mux_en_mscbus[2] = 1'b0;

assign DP1_3_in_mux_peripheral_mscbus[3] = io_SPI8CS3_out;

assign DP1_3_in_mux_en_mscbus[3] = io_SPI8CS3_oen;

// Assignments for DP1_3
assign io_SDFM1_i_datain1 = DP1_3_out_demux_peripheral_mscbus[1];

// Assignments for DP1_30
assign DP1_30_in_mux_peripheral_mscbus[1] = io_EPWM15_a_o;

assign DP1_30_in_mux_en_mscbus[1] = io_EPWM15_a_oen;

assign DP1_30_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR14_intr;

assign DP1_30_in_mux_en_mscbus[2] = 1'b0;

assign DP1_30_in_mux_peripheral_mscbus[4] = io_SPI3PICO_out;

assign DP1_30_in_mux_en_mscbus[4] = io_SPI3PICO_oen;

// Assignments for DP1_30
// Assignments for DP1_31
assign DP1_31_in_mux_peripheral_mscbus[1] = io_EPWM15_b_o;

assign DP1_31_in_mux_en_mscbus[1] = io_EPWM15_b_oen;

assign DP1_31_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR15_intr;

assign DP1_31_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_31
assign io_SPI3POCI_in = DP1_31_out_demux_peripheral_mscbus[1];

// Assignments for DP1_4
assign DP1_4_in_mux_peripheral_mscbus[1] = io_EPWM2_a_o;

assign DP1_4_in_mux_en_mscbus[1] = io_EPWM2_a_oen;

assign DP1_4_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR4_intr;

assign DP1_4_in_mux_en_mscbus[2] = 1'b0;

assign DP1_4_in_mux_peripheral_mscbus[3] = io_SPI8CLK_clock;

assign DP1_4_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP1_4
assign io_SDFM2_i_clock1 = DP1_4_out_demux_peripheral_mscbus[1];

// Assignments for DP1_5
assign DP1_5_in_mux_peripheral_mscbus[1] = io_EPWM2_b_o;

assign DP1_5_in_mux_en_mscbus[1] = io_EPWM2_b_oen;

assign DP1_5_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR5_intr;

assign DP1_5_in_mux_en_mscbus[2] = 1'b0;

assign DP1_5_in_mux_peripheral_mscbus[3] = io_SPI8PICO_out;

assign DP1_5_in_mux_en_mscbus[3] = io_SPI8PICO_oen;

// Assignments for DP1_5
assign io_SDFM2_i_datain1 = DP1_5_out_demux_peripheral_mscbus[1];

// Assignments for DP1_6
assign DP1_6_in_mux_peripheral_mscbus[1] = io_EPWM3_a_o;

assign DP1_6_in_mux_en_mscbus[1] = io_EPWM3_a_oen;

assign DP1_6_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR6_intr;

assign DP1_6_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP1_6
assign io_SDFM3_i_clock1 = DP1_6_out_demux_peripheral_mscbus[1];

assign io_SPI8POCI_in = DP1_6_out_demux_peripheral_mscbus[2];

// Assignments for DP1_7
assign DP1_7_in_mux_peripheral_mscbus[1] = io_EPWM3_b_o;

assign DP1_7_in_mux_en_mscbus[1] = io_EPWM3_b_oen;

assign DP1_7_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR7_intr;

assign DP1_7_in_mux_en_mscbus[2] = 1'b0;

assign DP1_7_in_mux_peripheral_mscbus[3] = io_SPI8CS0_out;

assign DP1_7_in_mux_en_mscbus[3] = io_SPI8CS0_oen;

// Assignments for DP1_7
assign io_SDFM3_i_datain1 = DP1_7_out_demux_peripheral_mscbus[1];

// Assignments for DP1_8
assign DP1_8_in_mux_peripheral_mscbus[1] = io_EPWM4_a_o;

assign DP1_8_in_mux_en_mscbus[1] = io_EPWM4_a_oen;

assign DP1_8_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR8_intr;

assign DP1_8_in_mux_en_mscbus[2] = 1'b0;

assign DP1_8_in_mux_peripheral_mscbus[3] = io_SPI8CS1_out;

assign DP1_8_in_mux_en_mscbus[3] = io_SPI8CS1_oen;

// Assignments for DP1_8
assign io_SDFM4_i_clock1 = DP1_8_out_demux_peripheral_mscbus[1];

// Assignments for DP1_9
assign DP1_9_in_mux_peripheral_mscbus[1] = io_EPWM4_b_o;

assign DP1_9_in_mux_en_mscbus[1] = io_EPWM4_b_oen;

assign DP1_9_in_mux_peripheral_mscbus[2] = io_OUTPUTXBAR9_intr;

assign DP1_9_in_mux_en_mscbus[2] = 1'b0;

assign DP1_9_in_mux_peripheral_mscbus[3] = io_SPI8CS2_out;

assign DP1_9_in_mux_en_mscbus[3] = io_SPI8CS2_oen;

// Assignments for DP1_9
assign io_SDFM4_i_datain1 = DP1_9_out_demux_peripheral_mscbus[1];

// Assignments for DP2_0
assign DP2_0_in_mux_peripheral_mscbus[1] = io_EPWM16_a_o;

assign DP2_0_in_mux_en_mscbus[1] = io_EPWM16_a_oen;

assign DP2_0_in_mux_peripheral_mscbus[4] = io_SPI3CS0_out;

assign DP2_0_in_mux_en_mscbus[4] = io_SPI3CS0_oen;

// Assignments for DP2_0
// Assignments for DP2_1
assign DP2_1_in_mux_peripheral_mscbus[1] = io_EPWM16_b_o;

assign DP2_1_in_mux_en_mscbus[1] = io_EPWM16_b_oen;

assign DP2_1_in_mux_peripheral_mscbus[4] = io_SPI3CS1_out;

assign DP2_1_in_mux_en_mscbus[4] = io_SPI3CS1_oen;

// Assignments for DP2_1
// Assignments for DP2_10
assign DP2_10_in_mux_peripheral_mscbus[1] = io_EPWM21_a_o;

assign DP2_10_in_mux_en_mscbus[1] = io_EPWM21_a_oen;

assign DP2_10_in_mux_peripheral_mscbus[4] = io_SPI4CS3_out;

assign DP2_10_in_mux_en_mscbus[4] = io_SPI4CS3_oen;

// Assignments for DP2_10
// Assignments for DP2_11
assign DP2_11_in_mux_peripheral_mscbus[1] = io_EPWM21_b_o;

assign DP2_11_in_mux_en_mscbus[1] = io_EPWM21_b_oen;

assign DP2_11_in_mux_peripheral_mscbus[3] = io_SPI5CLK_clock;

assign DP2_11_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP2_11
// Assignments for DP2_12
assign DP2_12_in_mux_peripheral_mscbus[1] = io_EPWM22_a_o;

assign DP2_12_in_mux_en_mscbus[1] = io_EPWM22_a_oen;

assign DP2_12_in_mux_peripheral_mscbus[3] = io_SPI5PICO_out;

assign DP2_12_in_mux_en_mscbus[3] = io_SPI5PICO_oen;

assign DP2_12_in_mux_peripheral_mscbus[4] = io_FSI1TX_ck;

assign DP2_12_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP2_12
// Assignments for DP2_13
assign DP2_13_in_mux_peripheral_mscbus[1] = io_EPWM22_b_o;

assign DP2_13_in_mux_en_mscbus[1] = io_EPWM22_b_oen;

assign DP2_13_in_mux_peripheral_mscbus[5] = io_FSI1TX_d0;

assign DP2_13_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP2_13
assign io_SPI5POCI_in = DP2_13_out_demux_peripheral_mscbus[2];

// Assignments for DP2_14
assign DP2_14_in_mux_peripheral_mscbus[1] = io_EPWM23_a_o;

assign DP2_14_in_mux_en_mscbus[1] = io_EPWM23_a_oen;

assign DP2_14_in_mux_peripheral_mscbus[4] = io_SPI5CS0_out;

assign DP2_14_in_mux_en_mscbus[4] = io_SPI5CS0_oen;

assign DP2_14_in_mux_peripheral_mscbus[6] = io_FSI1TX_d1;

assign DP2_14_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP2_14
// Assignments for DP2_15
assign DP2_15_in_mux_peripheral_mscbus[1] = io_EPWM23_b_o;

assign DP2_15_in_mux_en_mscbus[1] = io_EPWM23_b_oen;

assign DP2_15_in_mux_peripheral_mscbus[4] = io_SPI5CS1_out;

assign DP2_15_in_mux_en_mscbus[4] = io_SPI5CS1_oen;

// Assignments for DP2_15
assign io_FSI1RX_ck = DP2_15_out_demux_peripheral_mscbus[3];

// Assignments for DP2_16
assign DP2_16_in_mux_peripheral_mscbus[1] = io_EPWM24_a_o;

assign DP2_16_in_mux_en_mscbus[1] = io_EPWM24_a_oen;

assign DP2_16_in_mux_peripheral_mscbus[4] = io_SPI5CS2_out;

assign DP2_16_in_mux_en_mscbus[4] = io_SPI5CS2_oen;

// Assignments for DP2_16
assign io_FSI1RX_d0 = DP2_16_out_demux_peripheral_mscbus[3];

// Assignments for DP2_17
assign DP2_17_in_mux_peripheral_mscbus[1] = io_EPWM24_b_o;

assign DP2_17_in_mux_en_mscbus[1] = io_EPWM24_b_oen;

assign DP2_17_in_mux_peripheral_mscbus[4] = io_SPI5CS3_out;

assign DP2_17_in_mux_en_mscbus[4] = io_SPI5CS3_oen;

// Assignments for DP2_17
assign io_FSI1RX_d1 = DP2_17_out_demux_peripheral_mscbus[3];

// Assignments for DP2_18
assign DP2_18_in_mux_peripheral_mscbus[1] = io_EPWM25_a_o;

assign DP2_18_in_mux_en_mscbus[1] = io_EPWM25_a_oen;

assign DP2_18_in_mux_peripheral_mscbus[4] = io_SPI6CLK_clock;

assign DP2_18_in_mux_en_mscbus[4] = 1'b0;

assign DP2_18_in_mux_peripheral_mscbus[6] = io_FSI2TX_ck;

assign DP2_18_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP2_18
// Assignments for DP2_19
assign DP2_19_in_mux_peripheral_mscbus[1] = io_EPWM25_b_o;

assign DP2_19_in_mux_en_mscbus[1] = io_EPWM25_b_oen;

assign DP2_19_in_mux_peripheral_mscbus[4] = io_SPI6PICO_out;

assign DP2_19_in_mux_en_mscbus[4] = io_SPI6PICO_oen;

assign DP2_19_in_mux_peripheral_mscbus[6] = io_FSI2TX_d0;

assign DP2_19_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP2_19
// Assignments for DP2_2
assign DP2_2_in_mux_peripheral_mscbus[1] = io_EPWM17_a_o;

assign DP2_2_in_mux_en_mscbus[1] = io_EPWM17_a_oen;

assign DP2_2_in_mux_peripheral_mscbus[4] = io_SPI3CS2_out;

assign DP2_2_in_mux_en_mscbus[4] = io_SPI3CS2_oen;

// Assignments for DP2_2
// Assignments for DP2_20
assign DP2_20_in_mux_peripheral_mscbus[1] = io_EPWM26_a_o;

assign DP2_20_in_mux_en_mscbus[1] = io_EPWM26_a_oen;

assign DP2_20_in_mux_peripheral_mscbus[5] = io_FSI2TX_d1;

assign DP2_20_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP2_20
assign io_SPI6POCI_in = DP2_20_out_demux_peripheral_mscbus[2];

// Assignments for DP2_21
assign DP2_21_in_mux_peripheral_mscbus[1] = io_EPWM26_b_o;

assign DP2_21_in_mux_en_mscbus[1] = io_EPWM26_b_oen;

assign DP2_21_in_mux_peripheral_mscbus[2] = io_CAN6_txd;

assign DP2_21_in_mux_en_mscbus[2] = 1'b0;

assign DP2_21_in_mux_peripheral_mscbus[4] = io_SPI6CS0_out;

assign DP2_21_in_mux_en_mscbus[4] = io_SPI6CS0_oen;

assign DP2_21_in_mux_peripheral_mscbus[5] = io_SPI8CS4_out;

assign DP2_21_in_mux_en_mscbus[5] = io_SPI8CS4_oen;

// Assignments for DP2_21
// Assignments for DP2_22
assign DP2_22_in_mux_peripheral_mscbus[1] = io_EPWM27_a_o;

assign DP2_22_in_mux_en_mscbus[1] = io_EPWM27_a_oen;

assign DP2_22_in_mux_peripheral_mscbus[3] = io_SPI6CS1_out;

assign DP2_22_in_mux_en_mscbus[3] = io_SPI6CS1_oen;

assign DP2_22_in_mux_peripheral_mscbus[4] = io_SPI8CS5_out;

assign DP2_22_in_mux_en_mscbus[4] = io_SPI8CS5_oen;

// Assignments for DP2_22
assign io_CAN6_rxd = DP2_22_out_demux_peripheral_mscbus[1];

// Assignments for DP2_23
assign DP2_23_in_mux_peripheral_mscbus[1] = io_EPWM27_b_o;

assign DP2_23_in_mux_en_mscbus[1] = io_EPWM27_b_oen;

assign DP2_23_in_mux_peripheral_mscbus[2] = io_CAN7_txd;

assign DP2_23_in_mux_en_mscbus[2] = 1'b0;

assign DP2_23_in_mux_peripheral_mscbus[4] = io_SPI6CS2_out;

assign DP2_23_in_mux_en_mscbus[4] = io_SPI6CS2_oen;

assign DP2_23_in_mux_peripheral_mscbus[5] = io_SPI3CS4_out;

assign DP2_23_in_mux_en_mscbus[5] = io_SPI3CS4_oen;

// Assignments for DP2_23
// Assignments for DP2_24
assign DP2_24_in_mux_peripheral_mscbus[1] = io_EPWM28_a_o;

assign DP2_24_in_mux_en_mscbus[1] = io_EPWM28_a_oen;

assign DP2_24_in_mux_peripheral_mscbus[3] = io_SPI6CS3_out;

assign DP2_24_in_mux_en_mscbus[3] = io_SPI6CS3_oen;

assign DP2_24_in_mux_peripheral_mscbus[4] = io_SPI3CS5_out;

assign DP2_24_in_mux_en_mscbus[4] = io_SPI3CS5_oen;

// Assignments for DP2_24
assign io_CAN7_rxd = DP2_24_out_demux_peripheral_mscbus[1];

// Assignments for DP2_25
assign DP2_25_in_mux_peripheral_mscbus[1] = io_EPWM28_b_o;

assign DP2_25_in_mux_en_mscbus[1] = io_EPWM28_b_oen;

assign DP2_25_in_mux_peripheral_mscbus[2] = io_CAN8_txd;

assign DP2_25_in_mux_en_mscbus[2] = 1'b0;

assign DP2_25_in_mux_peripheral_mscbus[4] = io_SPI7CLK_clock;

assign DP2_25_in_mux_en_mscbus[4] = 1'b0;

assign DP2_25_in_mux_peripheral_mscbus[5] = io_LIN6_txd;

assign DP2_25_in_mux_en_mscbus[5] = io_LIN6_tr_en;

// Assignments for DP2_25
// Assignments for DP2_26
assign DP2_26_in_mux_peripheral_mscbus[1] = io_EPWM29_a_o;

assign DP2_26_in_mux_en_mscbus[1] = io_EPWM29_a_oen;

assign DP2_26_in_mux_peripheral_mscbus[2] = io_SPI6CLK_clock;

assign DP2_26_in_mux_en_mscbus[2] = 1'b0;

assign DP2_26_in_mux_peripheral_mscbus[3] = io_SPI7PICO_out;

assign DP2_26_in_mux_en_mscbus[3] = io_SPI7PICO_oen;

// Assignments for DP2_26
assign io_CAN8_rxd = DP2_26_out_demux_peripheral_mscbus[1];

assign io_LIN6_rxd = DP2_26_out_demux_peripheral_mscbus[2];

// Assignments for DP2_27
assign DP2_27_in_mux_peripheral_mscbus[1] = io_EPWM29_b_o;

assign DP2_27_in_mux_en_mscbus[1] = io_EPWM29_b_oen;

assign DP2_27_in_mux_peripheral_mscbus[2] = io_CAN9_txd;

assign DP2_27_in_mux_en_mscbus[2] = 1'b0;

assign DP2_27_in_mux_peripheral_mscbus[3] = io_SPI6PICO_out;

assign DP2_27_in_mux_en_mscbus[3] = io_SPI6PICO_oen;

assign DP2_27_in_mux_peripheral_mscbus[4] = io_LIN7_txd;

assign DP2_27_in_mux_en_mscbus[4] = io_LIN7_tr_en;

// Assignments for DP2_27
assign io_SPI7POCI_in = DP2_27_out_demux_peripheral_mscbus[1];

// Assignments for DP2_28
assign DP2_28_in_mux_peripheral_mscbus[1] = io_EPWM30_a_o;

assign DP2_28_in_mux_en_mscbus[1] = io_EPWM30_a_oen;

assign DP2_28_in_mux_peripheral_mscbus[2] = io_SPI7CS0_out;

assign DP2_28_in_mux_en_mscbus[2] = io_SPI7CS0_oen;

// Assignments for DP2_28
assign io_CAN9_rxd = DP2_28_out_demux_peripheral_mscbus[1];

assign io_SPI6POCI_in = DP2_28_out_demux_peripheral_mscbus[2];

assign io_LIN7_rxd = DP2_28_out_demux_peripheral_mscbus[3];

// Assignments for DP2_29
assign DP2_29_in_mux_peripheral_mscbus[1] = io_EPWM30_b_o;

assign DP2_29_in_mux_en_mscbus[1] = io_EPWM30_b_oen;

assign DP2_29_in_mux_peripheral_mscbus[2] = io_CAN10_txd;

assign DP2_29_in_mux_en_mscbus[2] = 1'b0;

assign DP2_29_in_mux_peripheral_mscbus[3] = io_SPI6CS0_out;

assign DP2_29_in_mux_en_mscbus[3] = io_SPI6CS0_oen;

assign DP2_29_in_mux_peripheral_mscbus[4] = io_SPI7CS1_out;

assign DP2_29_in_mux_en_mscbus[4] = io_SPI7CS1_oen;

// Assignments for DP2_29
assign io_SDFM7_i_clock1 = DP2_29_out_demux_peripheral_mscbus[1];

// Assignments for DP2_3
assign DP2_3_in_mux_peripheral_mscbus[1] = io_EPWM17_b_o;

assign DP2_3_in_mux_en_mscbus[1] = io_EPWM17_b_oen;

assign DP2_3_in_mux_peripheral_mscbus[4] = io_SPI3CS3_out;

assign DP2_3_in_mux_en_mscbus[4] = io_SPI3CS3_oen;

// Assignments for DP2_3
// Assignments for DP2_30
assign DP2_30_in_mux_peripheral_mscbus[1] = io_EPWM31_a_o;

assign DP2_30_in_mux_en_mscbus[1] = io_EPWM31_a_oen;

assign DP2_30_in_mux_peripheral_mscbus[2] = io_SPI6CS1_out;

assign DP2_30_in_mux_en_mscbus[2] = io_SPI6CS1_oen;

assign DP2_30_in_mux_peripheral_mscbus[3] = io_SPI7CS2_out;

assign DP2_30_in_mux_en_mscbus[3] = io_SPI7CS2_oen;

// Assignments for DP2_30
assign io_CAN10_rxd = DP2_30_out_demux_peripheral_mscbus[1];

assign io_SDFM7_i_datain1 = DP2_30_out_demux_peripheral_mscbus[2];

// Assignments for DP2_31
assign DP2_31_in_mux_peripheral_mscbus[1] = io_EPWM31_b_o;

assign DP2_31_in_mux_en_mscbus[1] = io_EPWM31_b_oen;

assign DP2_31_in_mux_peripheral_mscbus[2] = io_CAN11_txd;

assign DP2_31_in_mux_en_mscbus[2] = 1'b0;

assign DP2_31_in_mux_peripheral_mscbus[3] = io_SPI6CS2_out;

assign DP2_31_in_mux_en_mscbus[3] = io_SPI6CS2_oen;

assign DP2_31_in_mux_peripheral_mscbus[4] = io_SPI7CS3_out;

assign DP2_31_in_mux_en_mscbus[4] = io_SPI7CS3_oen;

// Assignments for DP2_31
assign io_SDFM0_i_clock1 = DP2_31_out_demux_peripheral_mscbus[1];

// Assignments for DP2_4
assign DP2_4_in_mux_peripheral_mscbus[1] = io_EPWM18_a_o;

assign DP2_4_in_mux_en_mscbus[1] = io_EPWM18_a_oen;

assign DP2_4_in_mux_peripheral_mscbus[4] = io_SPI4CLK_clock;

assign DP2_4_in_mux_en_mscbus[4] = 1'b0;

// Assignments for DP2_4
// Assignments for DP2_5
assign DP2_5_in_mux_peripheral_mscbus[1] = io_EPWM18_b_o;

assign DP2_5_in_mux_en_mscbus[1] = io_EPWM18_b_oen;

assign DP2_5_in_mux_peripheral_mscbus[4] = io_SPI4PICO_out;

assign DP2_5_in_mux_en_mscbus[4] = io_SPI4PICO_oen;

// Assignments for DP2_5
// Assignments for DP2_6
assign DP2_6_in_mux_peripheral_mscbus[1] = io_EPWM19_a_o;

assign DP2_6_in_mux_en_mscbus[1] = io_EPWM19_a_oen;

// Assignments for DP2_6
assign io_SPI4POCI_in = DP2_6_out_demux_peripheral_mscbus[1];

// Assignments for DP2_7
assign DP2_7_in_mux_peripheral_mscbus[1] = io_EPWM19_b_o;

assign DP2_7_in_mux_en_mscbus[1] = io_EPWM19_b_oen;

assign DP2_7_in_mux_peripheral_mscbus[4] = io_SPI4CS0_out;

assign DP2_7_in_mux_en_mscbus[4] = io_SPI4CS0_oen;

// Assignments for DP2_7
// Assignments for DP2_8
assign DP2_8_in_mux_peripheral_mscbus[1] = io_EPWM20_a_o;

assign DP2_8_in_mux_en_mscbus[1] = io_EPWM20_a_oen;

assign DP2_8_in_mux_peripheral_mscbus[4] = io_SPI4CS1_out;

assign DP2_8_in_mux_en_mscbus[4] = io_SPI4CS1_oen;

// Assignments for DP2_8
// Assignments for DP2_9
assign DP2_9_in_mux_peripheral_mscbus[1] = io_EPWM20_b_o;

assign DP2_9_in_mux_en_mscbus[1] = io_EPWM20_b_oen;

assign DP2_9_in_mux_peripheral_mscbus[4] = io_SPI4CS2_out;

assign DP2_9_in_mux_en_mscbus[4] = io_SPI4CS2_oen;

// Assignments for DP2_9
// Assignments for DP3_0
assign DP3_0_in_mux_peripheral_mscbus[2] = io_SPI6CS3_out;

assign DP3_0_in_mux_en_mscbus[2] = io_SPI6CS3_oen;

assign DP3_0_in_mux_peripheral_mscbus[3] = io_SPI8CLK_clock;

assign DP3_0_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP3_0
assign io_CAN11_rxd = DP3_0_out_demux_peripheral_mscbus[1];

assign io_SDFM0_i_datain1 = DP3_0_out_demux_peripheral_mscbus[2];

// Assignments for DP3_1
assign DP3_1_in_mux_peripheral_mscbus[1] = io_EPWM16_a_o;

assign DP3_1_in_mux_en_mscbus[1] = io_EPWM16_a_oen;

assign DP3_1_in_mux_peripheral_mscbus[2] = io_FSI3TX_d0;

assign DP3_1_in_mux_en_mscbus[2] = 1'b0;

assign DP3_1_in_mux_peripheral_mscbus[3] = io_SPI4CLK_clock;

assign DP3_1_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP3_1
assign io_SENT2_rxd_i = DP3_1_out_demux_peripheral_mscbus[1];

assign io_SPI5POCI_in = DP3_1_out_demux_peripheral_mscbus[2];

// Assignments for DP3_10
assign DP3_10_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS3_out;

assign DP3_10_in_mux_en_mscbus[1] = io_MIBSPI0CS3_oen;

assign DP3_10_in_mux_peripheral_mscbus[2] = io_EPWM20_b_o;

assign DP3_10_in_mux_en_mscbus[2] = io_EPWM20_b_oen;

assign DP3_10_in_mux_peripheral_mscbus[3] = io_PSI5_2_tx;

assign DP3_10_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP3_10
assign io_SPI4POCI_in = DP3_10_out_demux_peripheral_mscbus[1];

assign io_FSI4RX_d0 = DP3_10_out_demux_peripheral_mscbus[2];

assign io_SPI5POCI_in = DP3_10_out_demux_peripheral_mscbus[3];

// Assignments for DP3_11
assign DP3_11_in_mux_peripheral_mscbus[1] = io_MIBSPI1CLK_clock;

assign DP3_11_in_mux_en_mscbus[1] = 1'b0;

assign DP3_11_in_mux_peripheral_mscbus[2] = io_SPI3CS5_out;

assign DP3_11_in_mux_en_mscbus[2] = io_SPI3CS5_oen;

assign DP3_11_in_mux_peripheral_mscbus[3] = io_EPWM21_a_o;

assign DP3_11_in_mux_en_mscbus[3] = io_EPWM21_a_oen;

assign DP3_11_in_mux_peripheral_mscbus[4] = io_SPI5CS0_out;

assign DP3_11_in_mux_en_mscbus[4] = io_SPI5CS0_oen;

// Assignments for DP3_11
assign io_FSI4RX_d1 = DP3_11_out_demux_peripheral_mscbus[1];

assign io_PSI5_2_rx = DP3_11_out_demux_peripheral_mscbus[2];

// Assignments for DP3_12
assign DP3_12_in_mux_peripheral_mscbus[1] = io_MIBSPI1PICO_out;

assign DP3_12_in_mux_en_mscbus[1] = io_MIBSPI1PICO_oen;

assign DP3_12_in_mux_peripheral_mscbus[3] = io_EPWM21_b_o;

assign DP3_12_in_mux_en_mscbus[3] = io_EPWM21_b_oen;

assign DP3_12_in_mux_peripheral_mscbus[4] = io_FSI5TX_ck;

assign DP3_12_in_mux_en_mscbus[4] = 1'b0;

assign DP3_12_in_mux_peripheral_mscbus[5] = io_SPI5CS1_out;

assign DP3_12_in_mux_en_mscbus[5] = io_SPI5CS1_oen;

assign DP3_12_in_mux_peripheral_mscbus[6] = io_PSI5_3_tx;

assign DP3_12_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP3_12
// Assignments for DP3_13
assign DP3_13_in_mux_peripheral_mscbus[2] = io_EPWM22_a_o;

assign DP3_13_in_mux_en_mscbus[2] = io_EPWM22_a_oen;

assign DP3_13_in_mux_peripheral_mscbus[3] = io_FSI5TX_d0;

assign DP3_13_in_mux_en_mscbus[3] = 1'b0;

assign DP3_13_in_mux_peripheral_mscbus[4] = io_SPI5CS2_out;

assign DP3_13_in_mux_en_mscbus[4] = io_SPI5CS2_oen;

// Assignments for DP3_13
assign io_MIBSPI1POCI_in = DP3_13_out_demux_peripheral_mscbus[1];

assign io_PSI5_3_rx = DP3_13_out_demux_peripheral_mscbus[2];

// Assignments for DP3_14
assign DP3_14_in_mux_peripheral_mscbus[1] = io_MIBSPI1CS0_out;

assign DP3_14_in_mux_en_mscbus[1] = io_MIBSPI1CS0_oen;

assign DP3_14_in_mux_peripheral_mscbus[3] = io_EPWM22_b_o;

assign DP3_14_in_mux_en_mscbus[3] = io_EPWM22_b_oen;

assign DP3_14_in_mux_peripheral_mscbus[4] = io_FSI5TX_d1;

assign DP3_14_in_mux_en_mscbus[4] = 1'b0;

assign DP3_14_in_mux_peripheral_mscbus[5] = io_SPI5CS3_out;

assign DP3_14_in_mux_en_mscbus[5] = io_SPI5CS3_oen;

assign DP3_14_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS4_out;

assign DP3_14_in_mux_en_mscbus[6] = io_MIBSPI1CS4_oen;

// Assignments for DP3_14
// Assignments for DP3_15
assign DP3_15_in_mux_peripheral_mscbus[1] = io_MIBSPI1CS1_out;

assign DP3_15_in_mux_en_mscbus[1] = io_MIBSPI1CS1_oen;

assign DP3_15_in_mux_peripheral_mscbus[2] = io_SPI4CS0_out;

assign DP3_15_in_mux_en_mscbus[2] = io_SPI4CS0_oen;

assign DP3_15_in_mux_peripheral_mscbus[3] = io_EPWM23_a_o;

assign DP3_15_in_mux_en_mscbus[3] = io_EPWM23_a_oen;

assign DP3_15_in_mux_peripheral_mscbus[4] = io_SPI6CLK_clock;

assign DP3_15_in_mux_en_mscbus[4] = 1'b0;

assign DP3_15_in_mux_peripheral_mscbus[5] = io_MIBSPI1CS5_out;

assign DP3_15_in_mux_en_mscbus[5] = io_MIBSPI1CS5_oen;

// Assignments for DP3_15
assign io_FSI5RX_ck = DP3_15_out_demux_peripheral_mscbus[1];

// Assignments for DP3_16
assign DP3_16_in_mux_peripheral_mscbus[1] = io_MIBSPI1CS2_out;

assign DP3_16_in_mux_en_mscbus[1] = io_MIBSPI1CS2_oen;

assign DP3_16_in_mux_peripheral_mscbus[2] = io_SPI4CS1_out;

assign DP3_16_in_mux_en_mscbus[2] = io_SPI4CS1_oen;

assign DP3_16_in_mux_peripheral_mscbus[3] = io_EPWM23_b_o;

assign DP3_16_in_mux_en_mscbus[3] = io_EPWM23_b_oen;

assign DP3_16_in_mux_peripheral_mscbus[4] = io_SPI6PICO_out;

assign DP3_16_in_mux_en_mscbus[4] = io_SPI6PICO_oen;

assign DP3_16_in_mux_peripheral_mscbus[5] = io_MIBSPI1CS6_out;

assign DP3_16_in_mux_en_mscbus[5] = io_MIBSPI1CS6_oen;

// Assignments for DP3_16
assign io_FSI5RX_d0 = DP3_16_out_demux_peripheral_mscbus[1];

// Assignments for DP3_17
assign DP3_17_in_mux_peripheral_mscbus[2] = io_SPI4CS2_out;

assign DP3_17_in_mux_en_mscbus[2] = io_SPI4CS2_oen;

assign DP3_17_in_mux_peripheral_mscbus[3] = io_EPWM24_a_o;

assign DP3_17_in_mux_en_mscbus[3] = io_EPWM24_a_oen;

assign DP3_17_in_mux_peripheral_mscbus[4] = io_MIBSPI1CS7_out;

assign DP3_17_in_mux_en_mscbus[4] = io_MIBSPI1CS7_oen;

// Assignments for DP3_17
assign io_FSI5RX_d1 = DP3_17_out_demux_peripheral_mscbus[1];

assign io_SPI6POCI_in = DP3_17_out_demux_peripheral_mscbus[2];

// Assignments for DP3_18
assign DP3_18_in_mux_peripheral_mscbus[2] = io_SPI4CS3_out;

assign DP3_18_in_mux_en_mscbus[2] = io_SPI4CS3_oen;

assign DP3_18_in_mux_peripheral_mscbus[3] = io_EPWM24_b_o;

assign DP3_18_in_mux_en_mscbus[3] = io_EPWM24_b_oen;

assign DP3_18_in_mux_peripheral_mscbus[5] = io_SPI6CS0_out;

assign DP3_18_in_mux_en_mscbus[5] = io_SPI6CS0_oen;

assign DP3_18_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS8_out;

assign DP3_18_in_mux_en_mscbus[6] = io_MIBSPI1CS8_oen;

// Assignments for DP3_18
// Assignments for DP3_19
assign DP3_19_in_mux_peripheral_mscbus[3] = io_EPWM25_a_o;

assign DP3_19_in_mux_en_mscbus[3] = io_EPWM25_a_oen;

assign DP3_19_in_mux_peripheral_mscbus[5] = io_SPI6CS1_out;

assign DP3_19_in_mux_en_mscbus[5] = io_SPI6CS1_oen;

assign DP3_19_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS9_out;

assign DP3_19_in_mux_en_mscbus[6] = io_MIBSPI1CS9_oen;

// Assignments for DP3_19
// Assignments for DP3_2
assign DP3_2_in_mux_peripheral_mscbus[1] = io_SPI5CS0_out;

assign DP3_2_in_mux_en_mscbus[1] = io_SPI5CS0_oen;

assign DP3_2_in_mux_peripheral_mscbus[2] = io_EPWM16_b_o;

assign DP3_2_in_mux_en_mscbus[2] = io_EPWM16_b_oen;

assign DP3_2_in_mux_peripheral_mscbus[3] = io_FSI3TX_d1;

assign DP3_2_in_mux_en_mscbus[3] = 1'b0;

assign DP3_2_in_mux_peripheral_mscbus[4] = io_SPI4PICO_out;

assign DP3_2_in_mux_en_mscbus[4] = io_SPI4PICO_oen;

// Assignments for DP3_2
assign io_SENT3_rxd_i = DP3_2_out_demux_peripheral_mscbus[1];

// Assignments for DP3_20
assign DP3_20_in_mux_peripheral_mscbus[3] = io_EPWM25_b_o;

assign DP3_20_in_mux_en_mscbus[3] = io_EPWM25_b_oen;

assign DP3_20_in_mux_peripheral_mscbus[5] = io_SPI6CS2_out;

assign DP3_20_in_mux_en_mscbus[5] = io_SPI6CS2_oen;

assign DP3_20_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS10_out;

assign DP3_20_in_mux_en_mscbus[6] = io_MIBSPI1CS10_oen;

// Assignments for DP3_20
// Assignments for DP3_21
assign DP3_21_in_mux_peripheral_mscbus[3] = io_EPWM26_a_o;

assign DP3_21_in_mux_en_mscbus[3] = io_EPWM26_a_oen;

assign DP3_21_in_mux_peripheral_mscbus[5] = io_SPI6CS3_out;

assign DP3_21_in_mux_en_mscbus[5] = io_SPI6CS3_oen;

assign DP3_21_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS11_out;

assign DP3_21_in_mux_en_mscbus[6] = io_MIBSPI1CS11_oen;

// Assignments for DP3_21
// Assignments for DP3_22
assign DP3_22_in_mux_peripheral_mscbus[3] = io_EPWM26_b_o;

assign DP3_22_in_mux_en_mscbus[3] = io_EPWM26_b_oen;

assign DP3_22_in_mux_peripheral_mscbus[5] = io_EPWM31_b_o;

assign DP3_22_in_mux_en_mscbus[5] = io_EPWM31_b_oen;

assign DP3_22_in_mux_peripheral_mscbus[6] = io_SPI3CLK_clock;

assign DP3_22_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP3_22
// Assignments for DP3_23
assign DP3_23_in_mux_peripheral_mscbus[2] = io_FSI5TX_ck;

assign DP3_23_in_mux_en_mscbus[2] = 1'b0;

assign DP3_23_in_mux_peripheral_mscbus[3] = io_EPWM27_a_o;

assign DP3_23_in_mux_en_mscbus[3] = io_EPWM27_a_oen;

assign DP3_23_in_mux_peripheral_mscbus[5] = io_EPWM31_a_o;

assign DP3_23_in_mux_en_mscbus[5] = io_EPWM31_a_oen;

assign DP3_23_in_mux_peripheral_mscbus[6] = io_SPI3PICO_out;

assign DP3_23_in_mux_en_mscbus[6] = io_SPI3PICO_oen;

// Assignments for DP3_23
// Assignments for DP3_24
assign DP3_24_in_mux_peripheral_mscbus[2] = io_FSI5TX_d0;

assign DP3_24_in_mux_en_mscbus[2] = 1'b0;

assign DP3_24_in_mux_peripheral_mscbus[3] = io_EPWM27_b_o;

assign DP3_24_in_mux_en_mscbus[3] = io_EPWM27_b_oen;

assign DP3_24_in_mux_peripheral_mscbus[5] = io_EPWM30_b_o;

assign DP3_24_in_mux_en_mscbus[5] = io_EPWM30_b_oen;

// Assignments for DP3_24
assign io_SPI3POCI_in = DP3_24_out_demux_peripheral_mscbus[1];

// Assignments for DP3_25
assign DP3_25_in_mux_peripheral_mscbus[2] = io_FSI5TX_d1;

assign DP3_25_in_mux_en_mscbus[2] = 1'b0;

assign DP3_25_in_mux_peripheral_mscbus[3] = io_EPWM28_a_o;

assign DP3_25_in_mux_en_mscbus[3] = io_EPWM28_a_oen;

assign DP3_25_in_mux_peripheral_mscbus[5] = io_EPWM30_a_o;

assign DP3_25_in_mux_en_mscbus[5] = io_EPWM30_a_oen;

assign DP3_25_in_mux_peripheral_mscbus[6] = io_SPI3CS0_out;

assign DP3_25_in_mux_en_mscbus[6] = io_SPI3CS0_oen;

// Assignments for DP3_25
// Assignments for DP3_26
assign DP3_26_in_mux_peripheral_mscbus[2] = io_EPWM28_b_o;

assign DP3_26_in_mux_en_mscbus[2] = io_EPWM28_b_oen;

assign DP3_26_in_mux_peripheral_mscbus[4] = io_EPWM29_b_o;

assign DP3_26_in_mux_en_mscbus[4] = io_EPWM29_b_oen;

assign DP3_26_in_mux_peripheral_mscbus[5] = io_SPI3CS1_out;

assign DP3_26_in_mux_en_mscbus[5] = io_SPI3CS1_oen;

// Assignments for DP3_26
assign io_FSI5RX_ck = DP3_26_out_demux_peripheral_mscbus[1];

// Assignments for DP3_27
assign DP3_27_in_mux_peripheral_mscbus[2] = io_EPWM29_a_o;

assign DP3_27_in_mux_en_mscbus[2] = io_EPWM29_a_oen;

assign DP3_27_in_mux_peripheral_mscbus[4] = io_SPI3CS2_out;

assign DP3_27_in_mux_en_mscbus[4] = io_SPI3CS2_oen;

// Assignments for DP3_27
assign io_FSI5RX_d0 = DP3_27_out_demux_peripheral_mscbus[1];

// Assignments for DP3_28
assign DP3_28_in_mux_peripheral_mscbus[2] = io_EPWM29_b_o;

assign DP3_28_in_mux_en_mscbus[2] = io_EPWM29_b_oen;

assign DP3_28_in_mux_peripheral_mscbus[4] = io_EPWM28_b_o;

assign DP3_28_in_mux_en_mscbus[4] = io_EPWM28_b_oen;

assign DP3_28_in_mux_peripheral_mscbus[5] = io_SPI3CS3_out;

assign DP3_28_in_mux_en_mscbus[5] = io_SPI3CS3_oen;

// Assignments for DP3_28
assign io_FSI5RX_d1 = DP3_28_out_demux_peripheral_mscbus[1];

// Assignments for DP3_29
assign DP3_29_in_mux_peripheral_mscbus[1] = io_MIBSPI1CS3_out;

assign DP3_29_in_mux_en_mscbus[1] = io_MIBSPI1CS3_oen;

assign DP3_29_in_mux_peripheral_mscbus[2] = io_SPI8CLK_clock;

assign DP3_29_in_mux_en_mscbus[2] = 1'b0;

assign DP3_29_in_mux_peripheral_mscbus[5] = io_EPWM28_a_o;

assign DP3_29_in_mux_en_mscbus[5] = io_EPWM28_a_oen;

// Assignments for DP3_29
// Assignments for DP3_3
assign DP3_3_in_mux_peripheral_mscbus[1] = io_SPI5CS1_out;

assign DP3_3_in_mux_en_mscbus[1] = io_SPI5CS1_oen;

assign DP3_3_in_mux_peripheral_mscbus[2] = io_EPWM17_a_o;

assign DP3_3_in_mux_en_mscbus[2] = io_EPWM17_a_oen;

// Assignments for DP3_3
assign io_SENT4_rxd_i = DP3_3_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_ck = DP3_3_out_demux_peripheral_mscbus[2];

assign io_SPI4POCI_in = DP3_3_out_demux_peripheral_mscbus[3];

// Assignments for DP3_30
assign DP3_30_in_mux_peripheral_mscbus[1] = io_PSI5_0_tx;

assign DP3_30_in_mux_en_mscbus[1] = 1'b0;

assign DP3_30_in_mux_peripheral_mscbus[2] = io_SPI8PICO_out;

assign DP3_30_in_mux_en_mscbus[2] = io_SPI8PICO_oen;

assign DP3_30_in_mux_peripheral_mscbus[5] = io_EPWM27_b_o;

assign DP3_30_in_mux_en_mscbus[5] = io_EPWM27_b_oen;

// Assignments for DP3_30
// Assignments for DP3_31
assign DP3_31_in_mux_peripheral_mscbus[3] = io_EPWM27_a_o;

assign DP3_31_in_mux_en_mscbus[3] = io_EPWM27_a_oen;

// Assignments for DP3_31
assign io_PSI5_0_rx = DP3_31_out_demux_peripheral_mscbus[1];

assign io_SPI8POCI_in = DP3_31_out_demux_peripheral_mscbus[2];

// Assignments for DP3_4
assign DP3_4_in_mux_peripheral_mscbus[1] = io_MIBSPI0CLK_clock;

assign DP3_4_in_mux_en_mscbus[1] = 1'b0;

assign DP3_4_in_mux_peripheral_mscbus[2] = io_SPI5CS2_out;

assign DP3_4_in_mux_en_mscbus[2] = io_SPI5CS2_oen;

assign DP3_4_in_mux_peripheral_mscbus[3] = io_EPWM17_b_o;

assign DP3_4_in_mux_en_mscbus[3] = io_EPWM17_b_oen;

assign DP3_4_in_mux_peripheral_mscbus[4] = io_SPI4CS0_out;

assign DP3_4_in_mux_en_mscbus[4] = io_SPI4CS0_oen;

// Assignments for DP3_4
assign io_FSI3RX_d0 = DP3_4_out_demux_peripheral_mscbus[1];

// Assignments for DP3_5
assign DP3_5_in_mux_peripheral_mscbus[1] = io_MIBSPI0PICO_out;

assign DP3_5_in_mux_en_mscbus[1] = io_MIBSPI0PICO_oen;

assign DP3_5_in_mux_peripheral_mscbus[2] = io_SPI5CS3_out;

assign DP3_5_in_mux_en_mscbus[2] = io_SPI5CS3_oen;

assign DP3_5_in_mux_peripheral_mscbus[3] = io_EPWM18_a_o;

assign DP3_5_in_mux_en_mscbus[3] = io_EPWM18_a_oen;

assign DP3_5_in_mux_peripheral_mscbus[4] = io_SPI4CS1_out;

assign DP3_5_in_mux_en_mscbus[4] = io_SPI4CS1_oen;

// Assignments for DP3_5
assign io_FSI3RX_d1 = DP3_5_out_demux_peripheral_mscbus[1];

// Assignments for DP3_6
assign DP3_6_in_mux_peripheral_mscbus[1] = io_SPI3CS4_out;

assign DP3_6_in_mux_en_mscbus[1] = io_SPI3CS4_oen;

assign DP3_6_in_mux_peripheral_mscbus[2] = io_EPWM18_b_o;

assign DP3_6_in_mux_en_mscbus[2] = io_EPWM18_b_oen;

assign DP3_6_in_mux_peripheral_mscbus[3] = io_FSI4TX_ck;

assign DP3_6_in_mux_en_mscbus[3] = 1'b0;

assign DP3_6_in_mux_peripheral_mscbus[4] = io_SPI4CS2_out;

assign DP3_6_in_mux_en_mscbus[4] = io_SPI4CS2_oen;

// Assignments for DP3_6
assign io_MIBSPI0POCI_in = DP3_6_out_demux_peripheral_mscbus[1];

// Assignments for DP3_7
assign DP3_7_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS0_out;

assign DP3_7_in_mux_en_mscbus[1] = io_MIBSPI0CS0_oen;

assign DP3_7_in_mux_peripheral_mscbus[2] = io_EPWM19_a_o;

assign DP3_7_in_mux_en_mscbus[2] = io_EPWM19_a_oen;

assign DP3_7_in_mux_peripheral_mscbus[3] = io_FSI4TX_d0;

assign DP3_7_in_mux_en_mscbus[3] = 1'b0;

assign DP3_7_in_mux_peripheral_mscbus[4] = io_SPI4CS3_out;

assign DP3_7_in_mux_en_mscbus[4] = io_SPI4CS3_oen;

// Assignments for DP3_7
// Assignments for DP3_8
assign DP3_8_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS1_out;

assign DP3_8_in_mux_en_mscbus[1] = io_MIBSPI0CS1_oen;

assign DP3_8_in_mux_peripheral_mscbus[2] = io_SPI4CLK_clock;

assign DP3_8_in_mux_en_mscbus[2] = 1'b0;

assign DP3_8_in_mux_peripheral_mscbus[3] = io_EPWM19_b_o;

assign DP3_8_in_mux_en_mscbus[3] = io_EPWM19_b_oen;

assign DP3_8_in_mux_peripheral_mscbus[4] = io_FSI4TX_d1;

assign DP3_8_in_mux_en_mscbus[4] = 1'b0;

assign DP3_8_in_mux_peripheral_mscbus[5] = io_SPI5CLK_clock;

assign DP3_8_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP3_8
// Assignments for DP3_9
assign DP3_9_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS2_out;

assign DP3_9_in_mux_en_mscbus[1] = io_MIBSPI0CS2_oen;

assign DP3_9_in_mux_peripheral_mscbus[2] = io_SPI4PICO_out;

assign DP3_9_in_mux_en_mscbus[2] = io_SPI4PICO_oen;

assign DP3_9_in_mux_peripheral_mscbus[3] = io_EPWM20_a_o;

assign DP3_9_in_mux_en_mscbus[3] = io_EPWM20_a_oen;

assign DP3_9_in_mux_peripheral_mscbus[4] = io_SPI5PICO_out;

assign DP3_9_in_mux_en_mscbus[4] = io_SPI5PICO_oen;

// Assignments for DP3_9
assign io_FSI4RX_ck = DP3_9_out_demux_peripheral_mscbus[1];

// Assignments for DP4_0
assign DP4_0_in_mux_peripheral_mscbus[1] = io_PSI5_1_tx;

assign DP4_0_in_mux_en_mscbus[1] = 1'b0;

assign DP4_0_in_mux_peripheral_mscbus[2] = io_SPI8CS0_out;

assign DP4_0_in_mux_en_mscbus[2] = io_SPI8CS0_oen;

assign DP4_0_in_mux_peripheral_mscbus[5] = io_EPWM26_b_o;

assign DP4_0_in_mux_en_mscbus[5] = io_EPWM26_b_oen;

// Assignments for DP4_0
// Assignments for DP4_1
assign DP4_1_in_mux_peripheral_mscbus[1] = io_SPI8CS1_out;

assign DP4_1_in_mux_en_mscbus[1] = io_SPI8CS1_oen;

assign DP4_1_in_mux_peripheral_mscbus[4] = io_EPWM26_a_o;

assign DP4_1_in_mux_en_mscbus[4] = io_EPWM26_a_oen;

// Assignments for DP4_1
assign io_PSI5_1_rx = DP4_1_out_demux_peripheral_mscbus[1];

// Assignments for DP4_10
assign DP4_10_in_mux_peripheral_mscbus[2] = io_PSI5_1_tx;

assign DP4_10_in_mux_en_mscbus[2] = 1'b0;

assign DP4_10_in_mux_peripheral_mscbus[5] = io_EPWM21_b_o;

assign DP4_10_in_mux_en_mscbus[5] = io_EPWM21_b_oen;

// Assignments for DP4_10
assign io_MIBSPI0POCI_in = DP4_10_out_demux_peripheral_mscbus[2];

// Assignments for DP4_11
assign DP4_11_in_mux_peripheral_mscbus[4] = io_EPWM21_a_o;

assign DP4_11_in_mux_en_mscbus[4] = io_EPWM21_a_oen;

assign DP4_11_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS0_out;

assign DP4_11_in_mux_en_mscbus[5] = io_MIBSPI0CS0_oen;

// Assignments for DP4_11
assign io_PSI5_1_rx = DP4_11_out_demux_peripheral_mscbus[1];

// Assignments for DP4_12
assign DP4_12_in_mux_peripheral_mscbus[1] = io_FSI4TX_ck;

assign DP4_12_in_mux_en_mscbus[1] = 1'b0;

assign DP4_12_in_mux_peripheral_mscbus[4] = io_EPWM20_b_o;

assign DP4_12_in_mux_en_mscbus[4] = io_EPWM20_b_oen;

assign DP4_12_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS1_out;

assign DP4_12_in_mux_en_mscbus[5] = io_MIBSPI0CS1_oen;

// Assignments for DP4_12
// Assignments for DP4_13
assign DP4_13_in_mux_peripheral_mscbus[1] = io_FSI4TX_d0;

assign DP4_13_in_mux_en_mscbus[1] = 1'b0;

assign DP4_13_in_mux_peripheral_mscbus[4] = io_EPWM20_a_o;

assign DP4_13_in_mux_en_mscbus[4] = io_EPWM20_a_oen;

assign DP4_13_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS2_out;

assign DP4_13_in_mux_en_mscbus[5] = io_MIBSPI0CS2_oen;

// Assignments for DP4_13
// Assignments for DP4_14
assign DP4_14_in_mux_peripheral_mscbus[1] = io_FSI4TX_d1;

assign DP4_14_in_mux_en_mscbus[1] = 1'b0;

assign DP4_14_in_mux_peripheral_mscbus[4] = io_EPWM19_b_o;

assign DP4_14_in_mux_en_mscbus[4] = io_EPWM19_b_oen;

assign DP4_14_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS3_out;

assign DP4_14_in_mux_en_mscbus[5] = io_MIBSPI0CS3_oen;

// Assignments for DP4_14
// Assignments for DP4_15
assign DP4_15_in_mux_peripheral_mscbus[3] = io_EPWM19_a_o;

assign DP4_15_in_mux_en_mscbus[3] = io_EPWM19_a_oen;

assign DP4_15_in_mux_peripheral_mscbus[4] = io_MIBSPI0CS4_out;

assign DP4_15_in_mux_en_mscbus[4] = io_MIBSPI0CS4_oen;

// Assignments for DP4_15
assign io_FSI4RX_ck = DP4_15_out_demux_peripheral_mscbus[2];

assign io_SENT0_rxd_i = DP4_15_out_demux_peripheral_mscbus[3];

// Assignments for DP4_16
assign DP4_16_in_mux_peripheral_mscbus[3] = io_EPWM18_b_o;

assign DP4_16_in_mux_en_mscbus[3] = io_EPWM18_b_oen;

assign DP4_16_in_mux_peripheral_mscbus[4] = io_MIBSPI0CS5_out;

assign DP4_16_in_mux_en_mscbus[4] = io_MIBSPI0CS5_oen;

// Assignments for DP4_16
assign io_FSI4RX_d0 = DP4_16_out_demux_peripheral_mscbus[2];

assign io_SENT1_rxd_i = DP4_16_out_demux_peripheral_mscbus[3];

// Assignments for DP4_17
assign DP4_17_in_mux_peripheral_mscbus[3] = io_EPWM18_a_o;

assign DP4_17_in_mux_en_mscbus[3] = io_EPWM18_a_oen;

assign DP4_17_in_mux_peripheral_mscbus[4] = io_MIBSPI0CS6_out;

assign DP4_17_in_mux_en_mscbus[4] = io_MIBSPI0CS6_oen;

// Assignments for DP4_17
assign io_FSI4RX_d1 = DP4_17_out_demux_peripheral_mscbus[2];

assign io_SENT2_rxd_i = DP4_17_out_demux_peripheral_mscbus[3];

// Assignments for DP4_18
assign DP4_18_in_mux_peripheral_mscbus[1] = io_SPI2CS4_out;

assign DP4_18_in_mux_en_mscbus[1] = io_SPI2CS4_oen;

assign DP4_18_in_mux_peripheral_mscbus[2] = io_EPWM17_b_o;

assign DP4_18_in_mux_en_mscbus[2] = io_EPWM17_b_oen;

// Assignments for DP4_18
// Assignments for DP4_19
assign DP4_19_in_mux_peripheral_mscbus[2] = io_SPI2CS5_out;

assign DP4_19_in_mux_en_mscbus[2] = io_SPI2CS5_oen;

assign DP4_19_in_mux_peripheral_mscbus[4] = io_EPWM17_a_o;

assign DP4_19_in_mux_en_mscbus[4] = io_EPWM17_a_oen;

// Assignments for DP4_19
// Assignments for DP4_2
assign DP4_2_in_mux_peripheral_mscbus[1] = io_SPI3CLK_clock;

assign DP4_2_in_mux_en_mscbus[1] = 1'b0;

assign DP4_2_in_mux_peripheral_mscbus[2] = io_SPI8CS2_out;

assign DP4_2_in_mux_en_mscbus[2] = io_SPI8CS2_oen;

assign DP4_2_in_mux_peripheral_mscbus[5] = io_EPWM25_b_o;

assign DP4_2_in_mux_en_mscbus[5] = io_EPWM25_b_oen;

// Assignments for DP4_2
// Assignments for DP4_20
assign DP4_20_in_mux_peripheral_mscbus[3] = io_EPWM30_a_o;

assign DP4_20_in_mux_en_mscbus[3] = io_EPWM30_a_oen;

assign DP4_20_in_mux_peripheral_mscbus[5] = io_EPWM16_b_o;

assign DP4_20_in_mux_en_mscbus[5] = io_EPWM16_b_oen;

assign DP4_20_in_mux_peripheral_mscbus[6] = io_MIBSPI1CLK_clock;

assign DP4_20_in_mux_en_mscbus[6] = 1'b0;

assign DP4_20_in_mux_peripheral_mscbus[7] = io_MIBSPI0CS7_out;

assign DP4_20_in_mux_en_mscbus[7] = io_MIBSPI0CS7_oen;

// Assignments for DP4_20
// Assignments for DP4_21
assign DP4_21_in_mux_peripheral_mscbus[3] = io_EPWM30_b_o;

assign DP4_21_in_mux_en_mscbus[3] = io_EPWM30_b_oen;

assign DP4_21_in_mux_peripheral_mscbus[5] = io_EPWM16_a_o;

assign DP4_21_in_mux_en_mscbus[5] = io_EPWM16_a_oen;

assign DP4_21_in_mux_peripheral_mscbus[6] = io_MIBSPI1PICO_out;

assign DP4_21_in_mux_en_mscbus[6] = io_MIBSPI1PICO_oen;

assign DP4_21_in_mux_peripheral_mscbus[7] = io_MIBSPI0CS8_out;

assign DP4_21_in_mux_en_mscbus[7] = io_MIBSPI0CS8_oen;

// Assignments for DP4_21
// Assignments for DP4_22
assign DP4_22_in_mux_peripheral_mscbus[3] = io_EPWM31_a_o;

assign DP4_22_in_mux_en_mscbus[3] = io_EPWM31_a_oen;

assign DP4_22_in_mux_peripheral_mscbus[5] = io_EPWM15_b_o;

assign DP4_22_in_mux_en_mscbus[5] = io_EPWM15_b_oen;

assign DP4_22_in_mux_peripheral_mscbus[6] = io_MIBSPI0CS9_out;

assign DP4_22_in_mux_en_mscbus[6] = io_MIBSPI0CS9_oen;

// Assignments for DP4_22
assign io_MIBSPI1POCI_in = DP4_22_out_demux_peripheral_mscbus[2];

// Assignments for DP4_23
assign DP4_23_in_mux_peripheral_mscbus[3] = io_EPWM31_b_o;

assign DP4_23_in_mux_en_mscbus[3] = io_EPWM31_b_oen;

assign DP4_23_in_mux_peripheral_mscbus[5] = io_EPWM15_a_o;

assign DP4_23_in_mux_en_mscbus[5] = io_EPWM15_a_oen;

assign DP4_23_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS0_out;

assign DP4_23_in_mux_en_mscbus[6] = io_MIBSPI1CS0_oen;

assign DP4_23_in_mux_peripheral_mscbus[7] = io_MIBSPI0CS10_out;

assign DP4_23_in_mux_en_mscbus[7] = io_MIBSPI0CS10_oen;

// Assignments for DP4_23
// Assignments for DP4_24
assign DP4_24_in_mux_peripheral_mscbus[2] = io_LIN4_txd;

assign DP4_24_in_mux_en_mscbus[2] = io_LIN4_tr_en;

assign DP4_24_in_mux_peripheral_mscbus[5] = io_EPWM14_b_o;

assign DP4_24_in_mux_en_mscbus[5] = io_EPWM14_b_oen;

assign DP4_24_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS1_out;

assign DP4_24_in_mux_en_mscbus[6] = io_MIBSPI1CS1_oen;

assign DP4_24_in_mux_peripheral_mscbus[7] = io_MIBSPI0CS11_out;

assign DP4_24_in_mux_en_mscbus[7] = io_MIBSPI0CS11_oen;

// Assignments for DP4_24
// Assignments for DP4_25
assign DP4_25_in_mux_peripheral_mscbus[2] = io_SPI2CS4_out;

assign DP4_25_in_mux_en_mscbus[2] = io_SPI2CS4_oen;

assign DP4_25_in_mux_peripheral_mscbus[4] = io_EPWM14_a_o;

assign DP4_25_in_mux_en_mscbus[4] = io_EPWM14_a_oen;

assign DP4_25_in_mux_peripheral_mscbus[5] = io_MIBSPI1CS2_out;

assign DP4_25_in_mux_en_mscbus[5] = io_MIBSPI1CS2_oen;

// Assignments for DP4_25
assign io_LIN4_rxd = DP4_25_out_demux_peripheral_mscbus[2];

// Assignments for DP4_26
assign DP4_26_in_mux_peripheral_mscbus[2] = io_LIN5_txd;

assign DP4_26_in_mux_en_mscbus[2] = io_LIN5_tr_en;

assign DP4_26_in_mux_peripheral_mscbus[5] = io_EPWM13_b_o;

assign DP4_26_in_mux_en_mscbus[5] = io_EPWM13_b_oen;

assign DP4_26_in_mux_peripheral_mscbus[6] = io_MIBSPI1CS3_out;

assign DP4_26_in_mux_en_mscbus[6] = io_MIBSPI1CS3_oen;

// Assignments for DP4_26
// Assignments for DP4_27
assign DP4_27_in_mux_peripheral_mscbus[4] = io_EPWM13_a_o;

assign DP4_27_in_mux_en_mscbus[4] = io_EPWM13_a_oen;

assign DP4_27_in_mux_peripheral_mscbus[5] = io_SPI2CS5_out;

assign DP4_27_in_mux_en_mscbus[5] = io_SPI2CS5_oen;

// Assignments for DP4_27
assign io_LIN5_rxd = DP4_27_out_demux_peripheral_mscbus[2];

// Assignments for DP4_28
assign DP4_28_in_mux_peripheral_mscbus[2] = io_LIN6_txd;

assign DP4_28_in_mux_en_mscbus[2] = io_LIN6_tr_en;

assign DP4_28_in_mux_peripheral_mscbus[4] = io_EPWM12_b_o;

assign DP4_28_in_mux_en_mscbus[4] = io_EPWM12_b_oen;

assign DP4_28_in_mux_peripheral_mscbus[5] = io_CAN0_txd;

assign DP4_28_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP4_28
// Assignments for DP4_29
assign DP4_29_in_mux_peripheral_mscbus[4] = io_EPWM12_a_o;

assign DP4_29_in_mux_en_mscbus[4] = io_EPWM12_a_oen;

// Assignments for DP4_29
assign io_LIN6_rxd = DP4_29_out_demux_peripheral_mscbus[2];

assign io_CAN0_rxd = DP4_29_out_demux_peripheral_mscbus[3];

// Assignments for DP4_3
assign DP4_3_in_mux_peripheral_mscbus[1] = io_SPI3PICO_out;

assign DP4_3_in_mux_en_mscbus[1] = io_SPI3PICO_oen;

assign DP4_3_in_mux_peripheral_mscbus[2] = io_SPI8CS3_out;

assign DP4_3_in_mux_en_mscbus[2] = io_SPI8CS3_oen;

assign DP4_3_in_mux_peripheral_mscbus[5] = io_EPWM25_a_o;

assign DP4_3_in_mux_en_mscbus[5] = io_EPWM25_a_oen;

// Assignments for DP4_3
// Assignments for DP4_30
assign DP4_30_in_mux_peripheral_mscbus[4] = io_EPWM11_b_o;

assign DP4_30_in_mux_en_mscbus[4] = io_EPWM11_b_oen;

assign DP4_30_in_mux_peripheral_mscbus[5] = io_CAN1_txd;

assign DP4_30_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP4_30
assign io_SENT5_rxd_i = DP4_30_out_demux_peripheral_mscbus[2];

// Assignments for DP4_31
assign DP4_31_in_mux_peripheral_mscbus[4] = io_EPWM11_a_o;

assign DP4_31_in_mux_en_mscbus[4] = io_EPWM11_a_oen;

// Assignments for DP4_31
assign io_CAN1_rxd = DP4_31_out_demux_peripheral_mscbus[3];

// Assignments for DP4_4
assign DP4_4_in_mux_peripheral_mscbus[3] = io_EPWM24_b_o;

assign DP4_4_in_mux_en_mscbus[3] = io_EPWM24_b_oen;

assign DP4_4_in_mux_peripheral_mscbus[4] = io_SPI2CS4_out;

assign DP4_4_in_mux_en_mscbus[4] = io_SPI2CS4_oen;

// Assignments for DP4_4
assign io_SPI3POCI_in = DP4_4_out_demux_peripheral_mscbus[1];

// Assignments for DP4_5
assign DP4_5_in_mux_peripheral_mscbus[1] = io_SPI3CS0_out;

assign DP4_5_in_mux_en_mscbus[1] = io_SPI3CS0_oen;

assign DP4_5_in_mux_peripheral_mscbus[2] = io_SPI3CS1_out;

assign DP4_5_in_mux_en_mscbus[2] = io_SPI3CS1_oen;

assign DP4_5_in_mux_peripheral_mscbus[4] = io_EPWM24_a_o;

assign DP4_5_in_mux_en_mscbus[4] = io_EPWM24_a_oen;

assign DP4_5_in_mux_peripheral_mscbus[5] = io_SPI2CS5_out;

assign DP4_5_in_mux_en_mscbus[5] = io_SPI2CS5_oen;

// Assignments for DP4_5
// Assignments for DP4_6
assign DP4_6_in_mux_peripheral_mscbus[2] = io_SPI3CS2_out;

assign DP4_6_in_mux_en_mscbus[2] = io_SPI3CS2_oen;

assign DP4_6_in_mux_peripheral_mscbus[4] = io_EPWM23_b_o;

assign DP4_6_in_mux_en_mscbus[4] = io_EPWM23_b_oen;

assign DP4_6_in_mux_peripheral_mscbus[5] = io_UART1_tx;

assign DP4_6_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP4_6
// Assignments for DP4_7
assign DP4_7_in_mux_peripheral_mscbus[2] = io_SPI3CS3_out;

assign DP4_7_in_mux_en_mscbus[2] = io_SPI3CS3_oen;

assign DP4_7_in_mux_peripheral_mscbus[5] = io_EPWM23_a_o;

assign DP4_7_in_mux_en_mscbus[5] = io_EPWM23_a_oen;

// Assignments for DP4_7
assign io_UART1_rx = DP4_7_out_demux_peripheral_mscbus[2];

// Assignments for DP4_8
assign DP4_8_in_mux_peripheral_mscbus[2] = io_PSI5_0_tx;

assign DP4_8_in_mux_en_mscbus[2] = 1'b0;

assign DP4_8_in_mux_peripheral_mscbus[5] = io_EPWM22_b_o;

assign DP4_8_in_mux_en_mscbus[5] = io_EPWM22_b_oen;

assign DP4_8_in_mux_peripheral_mscbus[6] = io_MIBSPI0CLK_clock;

assign DP4_8_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP4_8
// Assignments for DP4_9
assign DP4_9_in_mux_peripheral_mscbus[4] = io_EPWM22_a_o;

assign DP4_9_in_mux_en_mscbus[4] = io_EPWM22_a_oen;

assign DP4_9_in_mux_peripheral_mscbus[5] = io_MIBSPI0PICO_out;

assign DP4_9_in_mux_en_mscbus[5] = io_MIBSPI0PICO_oen;

// Assignments for DP4_9
assign io_PSI5_0_rx = DP4_9_out_demux_peripheral_mscbus[1];

// Assignments for DP5_0
assign DP5_0_in_mux_peripheral_mscbus[2] = io_MIBSPI0CS2_out;

assign DP5_0_in_mux_en_mscbus[2] = io_MIBSPI0CS2_oen;

assign DP5_0_in_mux_peripheral_mscbus[5] = io_EPWM10_b_o;

assign DP5_0_in_mux_en_mscbus[5] = io_EPWM10_b_oen;

assign DP5_0_in_mux_peripheral_mscbus[6] = io_PSI5_0_tx;

assign DP5_0_in_mux_en_mscbus[6] = 1'b0;

assign DP5_0_in_mux_peripheral_mscbus[7] = io_SPI4CLK_clock;

assign DP5_0_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP5_0
// Assignments for DP5_1
assign DP5_1_in_mux_peripheral_mscbus[2] = io_MIBSPI0CS3_out;

assign DP5_1_in_mux_en_mscbus[2] = io_MIBSPI0CS3_oen;

assign DP5_1_in_mux_peripheral_mscbus[5] = io_EPWM10_a_o;

assign DP5_1_in_mux_en_mscbus[5] = io_EPWM10_b_oen;

assign DP5_1_in_mux_peripheral_mscbus[6] = io_SPI4PICO_out;

assign DP5_1_in_mux_en_mscbus[6] = io_SPI4PICO_oen;

// Assignments for DP5_1
assign io_PSI5_0_rx = DP5_1_out_demux_peripheral_mscbus[2];

// Assignments for DP5_10
assign DP5_10_in_mux_peripheral_mscbus[1] = io_MIBSPI0PICO_out;

assign DP5_10_in_mux_en_mscbus[1] = io_MIBSPI0PICO_oen;

assign DP5_10_in_mux_peripheral_mscbus[3] = io_SPI2CS0_out;

assign DP5_10_in_mux_en_mscbus[3] = io_SPI2CS0_oen;

assign DP5_10_in_mux_peripheral_mscbus[4] = io_EPWM5_b_o;

assign DP5_10_in_mux_en_mscbus[4] = io_EPWM5_b_oen;

assign DP5_10_in_mux_peripheral_mscbus[5] = io_SPI6CS0_out;

assign DP5_10_in_mux_en_mscbus[5] = io_SPI6CS0_oen;

// Assignments for DP5_10
// Assignments for DP5_11
assign DP5_11_in_mux_peripheral_mscbus[2] = io_SPI2CS1_out;

assign DP5_11_in_mux_en_mscbus[2] = io_SPI2CS1_oen;

assign DP5_11_in_mux_peripheral_mscbus[3] = io_EPWM5_a_o;

assign DP5_11_in_mux_en_mscbus[3] = io_EPWM5_a_oen;

assign DP5_11_in_mux_peripheral_mscbus[4] = io_SPI6CS1_out;

assign DP5_11_in_mux_en_mscbus[4] = io_SPI6CS1_oen;

// Assignments for DP5_11
assign io_MIBSPI0POCI_in = DP5_11_out_demux_peripheral_mscbus[2];

// Assignments for DP5_12
assign DP5_12_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS0_out;

assign DP5_12_in_mux_en_mscbus[1] = io_MIBSPI0CS0_oen;

assign DP5_12_in_mux_peripheral_mscbus[3] = io_SPI2CS2_out;

assign DP5_12_in_mux_en_mscbus[3] = io_SPI2CS2_oen;

assign DP5_12_in_mux_peripheral_mscbus[4] = io_EPWM4_b_o;

assign DP5_12_in_mux_en_mscbus[4] = io_EPWM4_b_oen;

assign DP5_12_in_mux_peripheral_mscbus[5] = io_SPI6CS2_out;

assign DP5_12_in_mux_en_mscbus[5] = io_SPI6CS2_oen;

// Assignments for DP5_12
// Assignments for DP5_13
assign DP5_13_in_mux_peripheral_mscbus[1] = io_MIBSPI0CS1_out;

assign DP5_13_in_mux_en_mscbus[1] = io_MIBSPI0CS1_oen;

assign DP5_13_in_mux_peripheral_mscbus[3] = io_SPI2CS3_out;

assign DP5_13_in_mux_en_mscbus[3] = io_SPI2CS3_oen;

assign DP5_13_in_mux_peripheral_mscbus[4] = io_EPWM4_a_o;

assign DP5_13_in_mux_en_mscbus[4] = io_EPWM4_a_oen;

assign DP5_13_in_mux_peripheral_mscbus[5] = io_SPI6CS3_out;

assign DP5_13_in_mux_en_mscbus[5] = io_SPI6CS3_oen;

// Assignments for DP5_13
// Assignments for DP5_14
assign DP5_14_in_mux_peripheral_mscbus[2] = io_CAN0_txd;

assign DP5_14_in_mux_en_mscbus[2] = 1'b0;

assign DP5_14_in_mux_peripheral_mscbus[5] = io_EPWM3_b_o;

assign DP5_14_in_mux_en_mscbus[5] = io_EPWM3_b_oen;

assign DP5_14_in_mux_peripheral_mscbus[6] = io_SPI7CLK_clock;

assign DP5_14_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP5_14
// Assignments for DP5_15
assign DP5_15_in_mux_peripheral_mscbus[4] = io_EPWM3_a_o;

assign DP5_15_in_mux_en_mscbus[4] = io_EPWM3_a_oen;

assign DP5_15_in_mux_peripheral_mscbus[5] = io_SPI7PICO_out;

assign DP5_15_in_mux_en_mscbus[5] = io_SPI7PICO_oen;

// Assignments for DP5_15
assign io_CAN0_rxd = DP5_15_out_demux_peripheral_mscbus[1];

// Assignments for DP5_16
assign DP5_16_in_mux_peripheral_mscbus[2] = io_CAN1_txd;

assign DP5_16_in_mux_en_mscbus[2] = 1'b0;

assign DP5_16_in_mux_peripheral_mscbus[5] = io_EPWM2_b_o;

assign DP5_16_in_mux_en_mscbus[5] = io_EPWM2_b_oen;

// Assignments for DP5_16
assign io_SPI7POCI_in = DP5_16_out_demux_peripheral_mscbus[1];

// Assignments for DP5_17
assign DP5_17_in_mux_peripheral_mscbus[4] = io_EPWM2_a_o;

assign DP5_17_in_mux_en_mscbus[4] = io_EPWM2_a_oen;

assign DP5_17_in_mux_peripheral_mscbus[5] = io_SPI7CS0_out;

assign DP5_17_in_mux_en_mscbus[5] = io_SPI7CS0_oen;

// Assignments for DP5_17
assign io_CAN1_rxd = DP5_17_out_demux_peripheral_mscbus[1];

// Assignments for DP5_18
assign DP5_18_in_mux_peripheral_mscbus[2] = io_CAN2_txd;

assign DP5_18_in_mux_en_mscbus[2] = 1'b0;

assign DP5_18_in_mux_peripheral_mscbus[4] = io_EPWM1_b_o;

assign DP5_18_in_mux_en_mscbus[4] = io_EPWM1_a_oen;

assign DP5_18_in_mux_peripheral_mscbus[5] = io_SPI7CS1_out;

assign DP5_18_in_mux_en_mscbus[5] = io_SPI7CS1_oen;

// Assignments for DP5_18
// Assignments for DP5_19
assign DP5_19_in_mux_peripheral_mscbus[3] = io_EPWM1_a_o;

assign DP5_19_in_mux_en_mscbus[3] = io_EPWM1_a_oen;

assign DP5_19_in_mux_peripheral_mscbus[4] = io_SPI7CS2_out;

assign DP5_19_in_mux_en_mscbus[4] = io_SPI7CS2_oen;

// Assignments for DP5_19
assign io_CAN2_rxd = DP5_19_out_demux_peripheral_mscbus[1];

// Assignments for DP5_2
assign DP5_2_in_mux_peripheral_mscbus[2] = io_SPI9CLK_clock;

assign DP5_2_in_mux_en_mscbus[2] = 1'b0;

assign DP5_2_in_mux_peripheral_mscbus[4] = io_EPWM9_b_o;

assign DP5_2_in_mux_en_mscbus[4] = io_EPWM9_b_oen;

assign DP5_2_in_mux_peripheral_mscbus[5] = io_PSI5_1_tx;

assign DP5_2_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP5_2
assign io_SPI4POCI_in = DP5_2_out_demux_peripheral_mscbus[1];

// Assignments for DP5_20
assign DP5_20_in_mux_peripheral_mscbus[1] = io_SPI2CLK_clock;

assign DP5_20_in_mux_en_mscbus[1] = 1'b0;

assign DP5_20_in_mux_peripheral_mscbus[2] = io_CAN3_txd;

assign DP5_20_in_mux_en_mscbus[2] = 1'b0;

assign DP5_20_in_mux_peripheral_mscbus[5] = io_EPWM0_b_o;

assign DP5_20_in_mux_en_mscbus[5] = io_EPWM0_b_oen;

assign DP5_20_in_mux_peripheral_mscbus[6] = io_SPI7CS3_out;

assign DP5_20_in_mux_en_mscbus[6] = io_SPI7CS3_oen;

// Assignments for DP5_20
// Assignments for DP5_21
assign DP5_21_in_mux_peripheral_mscbus[1] = io_SPI2PICO_out;

assign DP5_21_in_mux_en_mscbus[1] = io_SPI2PICO_oen;

assign DP5_21_in_mux_peripheral_mscbus[4] = io_EPWM0_a_o;

assign DP5_21_in_mux_en_mscbus[4] = io_EPWM0_a_oen;

assign DP5_21_in_mux_peripheral_mscbus[5] = io_PSI5_3_tx;

assign DP5_21_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP5_21
assign io_CAN3_rxd = DP5_21_out_demux_peripheral_mscbus[1];

// Assignments for DP5_22
assign DP5_22_in_mux_peripheral_mscbus[1] = io_CAN4_txd;

assign DP5_22_in_mux_en_mscbus[1] = 1'b0;

assign DP5_22_in_mux_peripheral_mscbus[4] = io_EPWM0_a_o;

assign DP5_22_in_mux_en_mscbus[4] = io_EPWM0_a_oen;

// Assignments for DP5_22
assign io_SPI2POCI_in = DP5_22_out_demux_peripheral_mscbus[1];

assign io_PSI5_3_rx = DP5_22_out_demux_peripheral_mscbus[2];

// Assignments for DP5_23
assign DP5_23_in_mux_peripheral_mscbus[1] = io_SPI2CS0_out;

assign DP5_23_in_mux_en_mscbus[1] = io_SPI2CS0_oen;

assign DP5_23_in_mux_peripheral_mscbus[4] = io_PSI5_2_tx;

assign DP5_23_in_mux_en_mscbus[4] = 1'b0;

assign DP5_23_in_mux_peripheral_mscbus[5] = io_SPI5CS1_out;

assign DP5_23_in_mux_en_mscbus[5] = io_SPI5CS1_oen;

// Assignments for DP5_23
assign io_CAN4_rxd = DP5_23_out_demux_peripheral_mscbus[1];

// Assignments for DP5_24
assign DP5_24_in_mux_peripheral_mscbus[1] = io_CAN5_txd;

assign DP5_24_in_mux_en_mscbus[1] = 1'b0;

assign DP5_24_in_mux_peripheral_mscbus[2] = io_SPI2CS1_out;

assign DP5_24_in_mux_en_mscbus[2] = io_SPI2CS1_oen;

assign DP5_24_in_mux_peripheral_mscbus[5] = io_SPI5CS2_out;

assign DP5_24_in_mux_en_mscbus[5] = io_SPI5CS2_oen;

// Assignments for DP5_24
assign io_PSI5_2_rx = DP5_24_out_demux_peripheral_mscbus[1];

// Assignments for DP5_25
assign DP5_25_in_mux_peripheral_mscbus[1] = io_SPI2CS2_out;

assign DP5_25_in_mux_en_mscbus[1] = io_SPI2CS2_oen;

assign DP5_25_in_mux_peripheral_mscbus[4] = io_SPI5CS3_out;

assign DP5_25_in_mux_en_mscbus[4] = io_SPI5CS3_oen;

// Assignments for DP5_25
assign io_CAN5_rxd = DP5_25_out_demux_peripheral_mscbus[1];

// Assignments for DP5_26
assign DP5_26_in_mux_peripheral_mscbus[2] = io_SPI2CS3_out;

assign DP5_26_in_mux_en_mscbus[2] = io_SPI2CS3_oen;

assign DP5_26_in_mux_peripheral_mscbus[5] = io_MIBSPI1CLK_clock;

assign DP5_26_in_mux_en_mscbus[5] = 1'b0;

assign DP5_26_in_mux_peripheral_mscbus[6] = io_EPWM24_a_o;

assign DP5_26_in_mux_en_mscbus[6] = io_EPWM24_a_oen;

// Assignments for DP5_26
// Assignments for DP5_27
assign DP5_27_in_mux_peripheral_mscbus[2] = io_FSI1TX_ck;

assign DP5_27_in_mux_en_mscbus[2] = 1'b0;

assign DP5_27_in_mux_peripheral_mscbus[5] = io_MIBSPI1PICO_out;

assign DP5_27_in_mux_en_mscbus[5] = io_MIBSPI1PICO_oen;

assign DP5_27_in_mux_peripheral_mscbus[6] = io_EPWM24_b_o;

assign DP5_27_in_mux_en_mscbus[6] = io_EPWM24_b_oen;

assign DP5_27_in_mux_peripheral_mscbus[7] = io_PSI5_3_tx;

assign DP5_27_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP5_27
// Assignments for DP5_28
assign DP5_28_in_mux_peripheral_mscbus[2] = io_FSI1TX_d0;

assign DP5_28_in_mux_en_mscbus[2] = 1'b0;

assign DP5_28_in_mux_peripheral_mscbus[5] = io_EPWM25_a_o;

assign DP5_28_in_mux_en_mscbus[5] = io_EPWM25_a_oen;

// Assignments for DP5_28
assign io_MIBSPI1POCI_in = DP5_28_out_demux_peripheral_mscbus[1];

assign io_PSI5_3_rx = DP5_28_out_demux_peripheral_mscbus[2];

// Assignments for DP5_29
assign DP5_29_in_mux_peripheral_mscbus[2] = io_FSI1TX_d1;

assign DP5_29_in_mux_en_mscbus[2] = 1'b0;

assign DP5_29_in_mux_peripheral_mscbus[5] = io_MIBSPI1CS0_out;

assign DP5_29_in_mux_en_mscbus[5] = io_MIBSPI1CS0_oen;

assign DP5_29_in_mux_peripheral_mscbus[6] = io_EPWM25_b_o;

assign DP5_29_in_mux_en_mscbus[6] = io_EPWM25_b_oen;

assign DP5_29_in_mux_peripheral_mscbus[7] = io_PSI5_2_tx;

assign DP5_29_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP5_29
// Assignments for DP5_3
assign DP5_3_in_mux_peripheral_mscbus[2] = io_SPI9PICO_out;

assign DP5_3_in_mux_en_mscbus[2] = io_SPI9PICO_oen;

assign DP5_3_in_mux_peripheral_mscbus[4] = io_EPWM9_a_o;

assign DP5_3_in_mux_en_mscbus[4] = io_EPWM9_a_oen;

assign DP5_3_in_mux_peripheral_mscbus[5] = io_SPI4CS0_out;

assign DP5_3_in_mux_en_mscbus[5] = io_SPI4CS0_oen;

// Assignments for DP5_3
assign io_PSI5_1_rx = DP5_3_out_demux_peripheral_mscbus[1];

// Assignments for DP5_30
assign DP5_30_in_mux_peripheral_mscbus[4] = io_MIBSPI1CS1_out;

assign DP5_30_in_mux_en_mscbus[4] = io_MIBSPI1CS1_oen;

assign DP5_30_in_mux_peripheral_mscbus[5] = io_EPWM26_a_o;

assign DP5_30_in_mux_en_mscbus[5] = io_EPWM26_a_oen;

// Assignments for DP5_30
assign io_FSI1RX_ck = DP5_30_out_demux_peripheral_mscbus[1];

assign io_PSI5_2_rx = DP5_30_out_demux_peripheral_mscbus[2];

// Assignments for DP5_31
assign DP5_31_in_mux_peripheral_mscbus[4] = io_MIBSPI1CS2_out;

assign DP5_31_in_mux_en_mscbus[4] = io_MIBSPI1CS2_oen;

assign DP5_31_in_mux_peripheral_mscbus[5] = io_EPWM26_b_o;

assign DP5_31_in_mux_en_mscbus[5] = io_EPWM26_b_oen;

assign DP5_31_in_mux_peripheral_mscbus[6] = io_SPI9CLK_clock;

assign DP5_31_in_mux_en_mscbus[6] = 1'b0;

assign DP5_31_in_mux_peripheral_mscbus[7] = io_PSI5_2_tx;

assign DP5_31_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP5_31
assign io_FSI1RX_d0 = DP5_31_out_demux_peripheral_mscbus[1];

// Assignments for DP5_4
assign DP5_4_in_mux_peripheral_mscbus[3] = io_LIN7_txd;

assign DP5_4_in_mux_en_mscbus[3] = io_LIN7_tr_en;

assign DP5_4_in_mux_peripheral_mscbus[4] = io_EPWM8_b_o;

assign DP5_4_in_mux_en_mscbus[4] = io_EPWM8_b_oen;

assign DP5_4_in_mux_peripheral_mscbus[5] = io_SPI4CS1_out;

assign DP5_4_in_mux_en_mscbus[5] = io_SPI4CS1_oen;

// Assignments for DP5_4
assign io_SPI9POCI_in = DP5_4_out_demux_peripheral_mscbus[1];

assign io_SENT3_rxd_i = DP5_4_out_demux_peripheral_mscbus[2];

// Assignments for DP5_5
assign DP5_5_in_mux_peripheral_mscbus[2] = io_SPI9CS0_out;

assign DP5_5_in_mux_en_mscbus[2] = io_SPI9CS0_oen;

assign DP5_5_in_mux_peripheral_mscbus[4] = io_EPWM8_a_o;

assign DP5_5_in_mux_en_mscbus[4] = io_EPWM8_a_oen;

assign DP5_5_in_mux_peripheral_mscbus[5] = io_SPI4CS2_out;

assign DP5_5_in_mux_en_mscbus[5] = io_SPI4CS2_oen;

// Assignments for DP5_5
assign io_LIN7_rxd = DP5_5_out_demux_peripheral_mscbus[1];

assign io_SENT4_rxd_i = DP5_5_out_demux_peripheral_mscbus[2];

// Assignments for DP5_6
assign DP5_6_in_mux_peripheral_mscbus[2] = io_SPI9CS1_out;

assign DP5_6_in_mux_en_mscbus[2] = io_SPI9CS1_oen;

assign DP5_6_in_mux_peripheral_mscbus[4] = io_MIBSPI1CS3_out;

assign DP5_6_in_mux_en_mscbus[4] = io_MIBSPI1CS3_oen;

assign DP5_6_in_mux_peripheral_mscbus[5] = io_EPWM7_b_o;

assign DP5_6_in_mux_en_mscbus[5] = io_EPWM7_b_oen;

assign DP5_6_in_mux_peripheral_mscbus[6] = io_SPI4CS3_out;

assign DP5_6_in_mux_en_mscbus[6] = io_SPI4CS3_oen;

// Assignments for DP5_6
assign io_SENT5_rxd_i = DP5_6_out_demux_peripheral_mscbus[1];

// Assignments for DP5_7
assign DP5_7_in_mux_peripheral_mscbus[2] = io_SPI9CS2_out;

assign DP5_7_in_mux_en_mscbus[2] = io_SPI9CS2_oen;

assign DP5_7_in_mux_peripheral_mscbus[4] = io_SPI2CLK_clock;

assign DP5_7_in_mux_en_mscbus[4] = 1'b0;

assign DP5_7_in_mux_peripheral_mscbus[5] = io_EPWM7_a_o;

assign DP5_7_in_mux_en_mscbus[5] = io_EPWM7_a_oen;

assign DP5_7_in_mux_peripheral_mscbus[6] = io_SPI6CLK_clock;

assign DP5_7_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP5_7
// Assignments for DP5_8
assign DP5_8_in_mux_peripheral_mscbus[1] = io_SPI9CS3_out;

assign DP5_8_in_mux_en_mscbus[1] = io_SPI9CS3_oen;

assign DP5_8_in_mux_peripheral_mscbus[3] = io_SPI2PICO_out;

assign DP5_8_in_mux_en_mscbus[3] = io_SPI2PICO_oen;

assign DP5_8_in_mux_peripheral_mscbus[4] = io_EPWM6_b_o;

assign DP5_8_in_mux_en_mscbus[4] = io_EPWM6_b_oen;

assign DP5_8_in_mux_peripheral_mscbus[5] = io_SPI6PICO_out;

assign DP5_8_in_mux_en_mscbus[5] = io_SPI6PICO_oen;

// Assignments for DP5_8
// Assignments for DP5_9
assign DP5_9_in_mux_peripheral_mscbus[1] = io_MIBSPI0CLK_clock;

assign DP5_9_in_mux_en_mscbus[1] = 1'b0;

assign DP5_9_in_mux_peripheral_mscbus[3] = io_EPWM6_a_o;

assign DP5_9_in_mux_en_mscbus[3] = io_EPWM6_a_oen;

// Assignments for DP5_9
assign io_SPI2POCI_in = DP5_9_out_demux_peripheral_mscbus[2];

assign io_SPI6POCI_in = DP5_9_out_demux_peripheral_mscbus[3];

// Assignments for DP6_0
assign DP6_0_in_mux_peripheral_mscbus[3] = io_MIBSPI1CS3_out;

assign DP6_0_in_mux_en_mscbus[3] = io_MIBSPI1CS3_oen;

assign DP6_0_in_mux_peripheral_mscbus[4] = io_SPI5CLK_clock;

assign DP6_0_in_mux_en_mscbus[4] = 1'b0;

assign DP6_0_in_mux_peripheral_mscbus[5] = io_SPI9PICO_out;

assign DP6_0_in_mux_en_mscbus[5] = io_SPI9PICO_oen;

// Assignments for DP6_0
assign io_FSI1RX_d1 = DP6_0_out_demux_peripheral_mscbus[2];

assign io_PSI5_2_rx = DP6_0_out_demux_peripheral_mscbus[3];

// Assignments for DP6_1
assign DP6_1_in_mux_peripheral_mscbus[1] = io_FSI2TX_ck;

assign DP6_1_in_mux_en_mscbus[1] = 1'b0;

assign DP6_1_in_mux_peripheral_mscbus[4] = io_SPI5PICO_out;

assign DP6_1_in_mux_en_mscbus[4] = io_SPI5PICO_oen;

assign DP6_1_in_mux_peripheral_mscbus[5] = io_PSI5_3_tx;

assign DP6_1_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP6_1
assign io_SPI9POCI_in = DP6_1_out_demux_peripheral_mscbus[2];

// Assignments for DP6_10
assign DP6_10_in_mux_peripheral_mscbus[2] = io_FSI3TX_d0;

assign DP6_10_in_mux_en_mscbus[2] = 1'b0;

assign DP6_10_in_mux_peripheral_mscbus[5] = io_EPWM3_a_o;

assign DP6_10_in_mux_en_mscbus[5] = io_EPWM3_a_oen;

assign DP6_10_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR6_intr;

assign DP6_10_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP6_10
// Assignments for DP6_11
assign DP6_11_in_mux_peripheral_mscbus[2] = io_FSI3TX_d1;

assign DP6_11_in_mux_en_mscbus[2] = 1'b0;

assign DP6_11_in_mux_peripheral_mscbus[6] = io_EPWM3_b_o;

assign DP6_11_in_mux_en_mscbus[6] = io_EPWM3_b_oen;

assign DP6_11_in_mux_peripheral_mscbus[7] = io_OUTPUTXBAR7_intr;

assign DP6_11_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP6_11
// Assignments for DP6_12
assign DP6_12_in_mux_peripheral_mscbus[1] = io_CAN5_txd;

assign DP6_12_in_mux_en_mscbus[1] = 1'b0;

assign DP6_12_in_mux_peripheral_mscbus[5] = io_EPWM24_a_o;

assign DP6_12_in_mux_en_mscbus[5] = io_EPWM24_a_oen;

assign DP6_12_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR8_intr;

assign DP6_12_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP6_12
// Assignments for DP6_13
assign DP6_13_in_mux_peripheral_mscbus[4] = io_EPWM24_b_o;

assign DP6_13_in_mux_en_mscbus[4] = io_EPWM24_b_oen;

assign DP6_13_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR9_intr;

assign DP6_13_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP6_13
assign io_CAN5_rxd = DP6_13_out_demux_peripheral_mscbus[2];

// Assignments for DP6_14
assign DP6_14_in_mux_peripheral_mscbus[5] = io_EPWM25_a_o;

assign DP6_14_in_mux_en_mscbus[5] = io_EPWM25_a_oen;

assign DP6_14_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR10_intr;

assign DP6_14_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP6_14
// Assignments for DP6_15
assign DP6_15_in_mux_peripheral_mscbus[4] = io_EPWM25_b_o;

assign DP6_15_in_mux_en_mscbus[4] = io_EPWM25_b_oen;

assign DP6_15_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR11_intr;

assign DP6_15_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP6_15
// Assignments for DP6_16
assign DP6_16_in_mux_peripheral_mscbus[5] = io_EPWM26_a_o;

assign DP6_16_in_mux_en_mscbus[5] = io_EPWM26_a_oen;

assign DP6_16_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR12_intr;

assign DP6_16_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP6_16
// Assignments for DP6_17
assign DP6_17_in_mux_peripheral_mscbus[6] = io_EPWM26_b_o;

assign DP6_17_in_mux_en_mscbus[6] = io_EPWM26_b_oen;

assign DP6_17_in_mux_peripheral_mscbus[7] = io_OUTPUTXBAR13_intr;

assign DP6_17_in_mux_en_mscbus[7] = 1'b0;

// Assignments for DP6_17
// Assignments for DP6_18
assign DP6_18_in_mux_peripheral_mscbus[5] = io_CAN2_txd;

assign DP6_18_in_mux_en_mscbus[5] = 1'b0;

assign DP6_18_in_mux_peripheral_mscbus[6] = io_MIBSPI0CS4_out;

assign DP6_18_in_mux_en_mscbus[6] = io_MIBSPI0CS4_oen;

// Assignments for DP6_18
// Assignments for DP6_19
assign DP6_19_in_mux_peripheral_mscbus[4] = io_SPI3CLK_clock;

assign DP6_19_in_mux_en_mscbus[4] = 1'b0;

assign DP6_19_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS5_out;

assign DP6_19_in_mux_en_mscbus[5] = io_MIBSPI0CS5_oen;

// Assignments for DP6_19
assign io_CAN2_rxd = DP6_19_out_demux_peripheral_mscbus[2];

// Assignments for DP6_2
assign DP6_2_in_mux_peripheral_mscbus[1] = io_FSI2TX_d0;

assign DP6_2_in_mux_en_mscbus[1] = 1'b0;

assign DP6_2_in_mux_peripheral_mscbus[5] = io_SPI9CS0_out;

assign DP6_2_in_mux_en_mscbus[5] = io_SPI9CS0_oen;

// Assignments for DP6_2
assign io_SPI5POCI_in = DP6_2_out_demux_peripheral_mscbus[2];

assign io_PSI5_3_rx = DP6_2_out_demux_peripheral_mscbus[3];

// Assignments for DP6_20
assign DP6_20_in_mux_peripheral_mscbus[5] = io_SPI3PICO_out;

assign DP6_20_in_mux_en_mscbus[5] = io_SPI3PICO_oen;

assign DP6_20_in_mux_peripheral_mscbus[6] = io_CAN3_txd;

assign DP6_20_in_mux_en_mscbus[6] = 1'b0;

assign DP6_20_in_mux_peripheral_mscbus[7] = io_MIBSPI0CS6_out;

assign DP6_20_in_mux_en_mscbus[7] = io_MIBSPI0CS6_oen;

// Assignments for DP6_20
// Assignments for DP6_21
assign DP6_21_in_mux_peripheral_mscbus[4] = io_MIBSPI0CS7_out;

assign DP6_21_in_mux_en_mscbus[4] = io_MIBSPI0CS7_oen;

// Assignments for DP6_21
assign io_SPI3POCI_in = DP6_21_out_demux_peripheral_mscbus[2];

assign io_CAN3_rxd = DP6_21_out_demux_peripheral_mscbus[3];

// Assignments for DP6_22
assign DP6_22_in_mux_peripheral_mscbus[3] = io_SPI3CS0_out;

assign DP6_22_in_mux_en_mscbus[3] = io_SPI3CS0_oen;

assign DP6_22_in_mux_peripheral_mscbus[4] = io_CAN4_txd;

assign DP6_22_in_mux_en_mscbus[4] = 1'b0;

assign DP6_22_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS8_out;

assign DP6_22_in_mux_en_mscbus[5] = io_MIBSPI0CS8_oen;

// Assignments for DP6_22
// Assignments for DP6_23
assign DP6_23_in_mux_peripheral_mscbus[5] = io_SPI3CS1_out;

assign DP6_23_in_mux_en_mscbus[5] = io_SPI3CS1_oen;

assign DP6_23_in_mux_peripheral_mscbus[6] = io_MIBSPI0CS9_out;

assign DP6_23_in_mux_en_mscbus[6] = io_MIBSPI0CS9_oen;

// Assignments for DP6_23
assign io_CAN4_rxd = DP6_23_out_demux_peripheral_mscbus[1];

// Assignments for DP6_24
assign DP6_24_in_mux_peripheral_mscbus[4] = io_SPI3CS2_out;

assign DP6_24_in_mux_en_mscbus[4] = io_SPI3CS2_oen;

assign DP6_24_in_mux_peripheral_mscbus[5] = io_CAN5_txd;

assign DP6_24_in_mux_en_mscbus[5] = 1'b0;

assign DP6_24_in_mux_peripheral_mscbus[6] = io_MIBSPI0CS10_out;

assign DP6_24_in_mux_en_mscbus[6] = io_MIBSPI0CS10_oen;

// Assignments for DP6_24
// Assignments for DP6_25
assign DP6_25_in_mux_peripheral_mscbus[4] = io_SPI3CS3_out;

assign DP6_25_in_mux_en_mscbus[4] = io_SPI3CS3_oen;

assign DP6_25_in_mux_peripheral_mscbus[5] = io_MIBSPI0CS11_out;

assign DP6_25_in_mux_en_mscbus[5] = io_MIBSPI0CS11_oen;

// Assignments for DP6_25
assign io_CAN5_rxd = DP6_25_out_demux_peripheral_mscbus[2];

// Assignments for DP6_26
// Assignments for DP6_26
// Assignments for DP6_27
// Assignments for DP6_27
// Assignments for DP6_3
assign DP6_3_in_mux_peripheral_mscbus[1] = io_FSI2TX_d1;

assign DP6_3_in_mux_en_mscbus[1] = 1'b0;

assign DP6_3_in_mux_peripheral_mscbus[5] = io_SPI5CS0_out;

assign DP6_3_in_mux_en_mscbus[5] = io_SPI5CS0_oen;

assign DP6_3_in_mux_peripheral_mscbus[6] = io_SPI9CS1_out;

assign DP6_3_in_mux_en_mscbus[6] = io_SPI9CS1_oen;

// Assignments for DP6_3
// Assignments for DP6_4
assign DP6_4_in_mux_peripheral_mscbus[5] = io_SPI9CS2_out;

assign DP6_4_in_mux_en_mscbus[5] = io_SPI9CS2_oen;

// Assignments for DP6_4
// Assignments for DP6_5
assign DP6_5_in_mux_peripheral_mscbus[5] = io_SPI9CS3_out;

assign DP6_5_in_mux_en_mscbus[5] = io_SPI9CS3_oen;

// Assignments for DP6_5
// Assignments for DP6_6
assign DP6_6_in_mux_peripheral_mscbus[5] = io_EPWM1_a_o;

assign DP6_6_in_mux_en_mscbus[5] = io_EPWM1_a_oen;

assign DP6_6_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR2_intr;

assign DP6_6_in_mux_en_mscbus[6] = 1'b0;

assign DP6_6_in_mux_peripheral_mscbus[7] = io_SPI9CS4_out;

assign DP6_6_in_mux_en_mscbus[7] = io_SPI9CS4_oen;

// Assignments for DP6_6
assign io_FSI2RX_ck = DP6_6_out_demux_peripheral_mscbus[2];

// Assignments for DP6_7
assign DP6_7_in_mux_peripheral_mscbus[5] = io_EPWM1_b_o;

assign DP6_7_in_mux_en_mscbus[5] = io_EPWM1_a_oen;

assign DP6_7_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR3_intr;

assign DP6_7_in_mux_en_mscbus[6] = 1'b0;

assign DP6_7_in_mux_peripheral_mscbus[7] = io_SPI9CS5_out;

assign DP6_7_in_mux_en_mscbus[7] = io_SPI9CS5_oen;

// Assignments for DP6_7
assign io_FSI2RX_d0 = DP6_7_out_demux_peripheral_mscbus[2];

// Assignments for DP6_8
assign DP6_8_in_mux_peripheral_mscbus[4] = io_EPWM2_a_o;

assign DP6_8_in_mux_en_mscbus[4] = io_EPWM2_a_oen;

assign DP6_8_in_mux_peripheral_mscbus[5] = io_OUTPUTXBAR4_intr;

assign DP6_8_in_mux_en_mscbus[5] = 1'b0;

// Assignments for DP6_8
assign io_FSI2RX_d1 = DP6_8_out_demux_peripheral_mscbus[2];

// Assignments for DP6_9
assign DP6_9_in_mux_peripheral_mscbus[2] = io_FSI3TX_ck;

assign DP6_9_in_mux_en_mscbus[2] = 1'b0;

assign DP6_9_in_mux_peripheral_mscbus[5] = io_EPWM2_b_o;

assign DP6_9_in_mux_en_mscbus[5] = io_EPWM2_b_oen;

assign DP6_9_in_mux_peripheral_mscbus[6] = io_OUTPUTXBAR5_intr;

assign DP6_9_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP6_9
// Assignments for DP7_0
assign DP7_0_in_mux_peripheral_mscbus[5] = io_SPI2CS4_out;

assign DP7_0_in_mux_en_mscbus[5] = io_SPI2CS4_oen;

assign DP7_0_in_mux_peripheral_mscbus[6] = io_SPI6CS4_out;

assign DP7_0_in_mux_en_mscbus[6] = io_SPI6CS4_oen;

// Assignments for DP7_0
// Assignments for DP7_1
assign DP7_1_in_mux_peripheral_mscbus[3] = io_SPI2CS5_out;

assign DP7_1_in_mux_en_mscbus[3] = io_SPI2CS5_oen;

assign DP7_1_in_mux_peripheral_mscbus[4] = io_SPI6CS5_out;

assign DP7_1_in_mux_en_mscbus[4] = io_SPI6CS5_oen;

// Assignments for DP7_1
// Assignments for DP7_10
// Assignments for DP7_10
assign io_SDFM8_i_clock1 = DP7_10_out_demux_peripheral_mscbus[1];

assign io_PSI5_0_rx = DP7_10_out_demux_peripheral_mscbus[2];

assign io_PSI5_1_rx = DP7_10_out_demux_peripheral_mscbus[3];

// Assignments for DP7_11
assign DP7_11_in_mux_peripheral_mscbus[1] = io_SPI8CS4_out;

assign DP7_11_in_mux_en_mscbus[1] = io_SPI8CS4_oen;

assign DP7_11_in_mux_peripheral_mscbus[3] = io_CAN9_txd;

assign DP7_11_in_mux_en_mscbus[3] = 1'b0;

// Assignments for DP7_11
assign io_SDFM8_i_datain1 = DP7_11_out_demux_peripheral_mscbus[1];

// Assignments for DP7_12
assign DP7_12_in_mux_peripheral_mscbus[1] = io_SPI8CS5_out;

assign DP7_12_in_mux_en_mscbus[1] = io_SPI8CS5_oen;

// Assignments for DP7_12
assign io_SDFM9_i_clock1 = DP7_12_out_demux_peripheral_mscbus[1];

assign io_CAN9_rxd = DP7_12_out_demux_peripheral_mscbus[2];

// Assignments for DP7_13
assign DP7_13_in_mux_peripheral_mscbus[2] = io_CAN10_txd;

assign DP7_13_in_mux_en_mscbus[2] = 1'b0;

// Assignments for DP7_13
assign io_SDFM9_i_datain1 = DP7_13_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_ck = DP7_13_out_demux_peripheral_mscbus[2];

// Assignments for DP7_14
// Assignments for DP7_14
assign io_SDFM10_i_clock1 = DP7_14_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_d0 = DP7_14_out_demux_peripheral_mscbus[2];

assign io_CAN10_rxd = DP7_14_out_demux_peripheral_mscbus[3];

// Assignments for DP7_15
// Assignments for DP7_15
assign io_SDFM10_i_datain1 = DP7_15_out_demux_peripheral_mscbus[1];

assign io_FSI3RX_d1 = DP7_15_out_demux_peripheral_mscbus[2];

// Assignments for DP7_2
assign DP7_2_in_mux_peripheral_mscbus[5] = io_EPWM21_a_o;

assign DP7_2_in_mux_en_mscbus[5] = io_EPWM21_a_oen;

assign DP7_2_in_mux_peripheral_mscbus[6] = io_SPI5CS4_out;

assign DP7_2_in_mux_en_mscbus[6] = io_SPI5CS4_oen;

// Assignments for DP7_2
// Assignments for DP7_3
assign DP7_3_in_mux_peripheral_mscbus[5] = io_EPWM21_b_o;

assign DP7_3_in_mux_en_mscbus[5] = io_EPWM21_b_oen;

assign DP7_3_in_mux_peripheral_mscbus[6] = io_SPI5CS5_out;

assign DP7_3_in_mux_en_mscbus[6] = io_SPI5CS5_oen;

// Assignments for DP7_3
// Assignments for DP7_4
assign DP7_4_in_mux_peripheral_mscbus[5] = io_EPWM22_a_o;

assign DP7_4_in_mux_en_mscbus[5] = io_EPWM22_a_oen;

assign DP7_4_in_mux_peripheral_mscbus[6] = io_SPI4CS4_out;

assign DP7_4_in_mux_en_mscbus[6] = io_SPI4CS4_oen;

// Assignments for DP7_4
// Assignments for DP7_5
assign DP7_5_in_mux_peripheral_mscbus[5] = io_EPWM22_b_o;

assign DP7_5_in_mux_en_mscbus[5] = io_EPWM22_b_oen;

assign DP7_5_in_mux_peripheral_mscbus[6] = io_SPI4CS5_out;

assign DP7_5_in_mux_en_mscbus[6] = io_SPI4CS5_oen;

// Assignments for DP7_5
// Assignments for DP7_6
assign DP7_6_in_mux_peripheral_mscbus[4] = io_EPWM23_a_o;

assign DP7_6_in_mux_en_mscbus[4] = io_EPWM23_a_oen;

assign DP7_6_in_mux_peripheral_mscbus[5] = io_SPI5CS4_out;

assign DP7_6_in_mux_en_mscbus[5] = io_SPI5CS4_oen;

// Assignments for DP7_6
// Assignments for DP7_7
assign DP7_7_in_mux_peripheral_mscbus[4] = io_EPWM23_b_o;

assign DP7_7_in_mux_en_mscbus[4] = io_EPWM23_b_oen;

assign DP7_7_in_mux_peripheral_mscbus[5] = io_SPI5CS5_out;

assign DP7_7_in_mux_en_mscbus[5] = io_SPI5CS5_oen;

// Assignments for DP7_7
// Assignments for DP7_8
assign DP7_8_in_mux_peripheral_mscbus[5] = io_EPWM24_a_o;

assign DP7_8_in_mux_en_mscbus[5] = io_EPWM24_a_oen;

// Assignments for DP7_8
// Assignments for DP7_9
assign DP7_9_in_mux_peripheral_mscbus[2] = io_PSI5_0_tx;

assign DP7_9_in_mux_en_mscbus[2] = 1'b0;

assign DP7_9_in_mux_peripheral_mscbus[4] = io_EPWM24_b_o;

assign DP7_9_in_mux_en_mscbus[4] = io_EPWM24_b_oen;

assign DP7_9_in_mux_peripheral_mscbus[6] = io_PSI5_1_tx;

assign DP7_9_in_mux_en_mscbus[6] = 1'b0;

// Assignments for DP7_9

endmodule


